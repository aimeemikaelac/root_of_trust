

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hO+5yTBv4yTuDa91Fg43q7XKSAwGklxmlANdmlwbT2i830ylPy5q/f79HNxzAKl6I+pBIq+6lJb6
Eg2EkCV5tA==


`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Fe8TkBtfpoMxA1zPCIfGNLiAp4jEfQh/goK0f75sgsYb8oM9g69RyvHQwgEF+/RM0w6/mzZ2TrlD
SHA2BSwfxzGGXZehRhmxFx0o3QsMeWKPS+wvqNpmxi9sig95TdAyIjQgccr++z/J1ffIQcnvgdgB
b8qacZ76DAzEAabXnxY=


`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
lAJ5QvJO/R06hMi30eQWGtinWISST/IjqTzxCGxltVzO7YNbbIYKonJJxaA8RjBMhwJZ2Pp3sTKe
Y3PPIPu8v0i4csjGysocsoLlymimxv1ZWNcI7QNgFS+BfRThzEf0tKuUU3FB92JF4E3vLuesYqBc
ydslg708Tme3kSkC7sY=


`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
qi6tHZ7LdgkxpjN1kl/XIM6fD7tPqvPdyItomOgwiMn8+LN+1Z7aaZt3+QF+cH0ZckOuf+LIqu/B
y+oF8DRJodEOj4k2FYG32dynnmByxOveiByRaqXl2TJBv+L1b3+qu5XaNndxDPIFdA1N6WkKbJyU
qW9QQrh6MAneTunUBnxPyKtf/vISgOenOHQH1BckT611EHdxIkF9XWrVL/xO6bdpWz37eKsxFcyI
SoO5/pXllalyNBWFkYuEzqwMM5YYlcO/EeTByldLQAoeGa4E9vxvz3Pnur3XC8dRL+wXI6tnaa3j
cGxWR77DWdQj+mUaLSw5JrUcQiX6kJDuRrwhmg==


`pragma protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
qO22OLKzHZSFCxUoDtULBmK+/f1CGSOef+wul05EHVTgo3G09WNIBDll00kfhmJkGec4DfrLQJsC
kN0k5vMZX0tHWgrX0EW2Ee1rAUZIF/fP2Fiivkj6xW3+hICMkvuZx9OGe2/XEYpvvZ+atbXIujgS
zrHx5LLRxvPVxsdY6y+8WhKT/xJQblT5FC6EEmvQcu6hW/gBloFIfKiFjUE7fI3ks4y9fdycSuMj
skuWheywhax+Cv+IloqibEl+LKiDgquLGUBCSrqkWweUaFGswNklrEAtVw0G6IgdB3YMO3M90edU
Na2OM57JX1nETEFj7JYWacF3yNpQ208t9MKy3w==


`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
oh34PooggCnD0DQrUODr3G1zyfO6UmERje/ryZcPsL6gFLTpWBHdkK0onoL141U9Wn3RBdoXSj1J
qL75oPfPY/R17F0ONnPnj/pxLgRXWaSgAEauOpU1uMuuS9mXIFqghCzCYn72U6M8a5QkbxwLjnzH
C1ks2XcXsRj2u3zIqAKykOqn/jPDDBOUSM4CS6ovKMy5VAszToUjI7pAScajaNXQg1gnvHC8lpTJ
4dI3+XNgFRx7Uh6JvDRJ/fFod0nFRpMUk4EPXxnpeoXC8FEcaZSJ2HQGAlzYacoxAXMwL0zLk1U6
oWqc0x7jViy9oDctKEUpdT8butOlm0XTDZfOeQ==


`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 568944)
`pragma protect data_block
ySTDCaxTcpQ6P79suOQEUzg/U+Ra59CytEXWfHm0NXQkNByNzw+I6XOpAnSvu/W1N/nhidlZ8De8
y/GNuI2YWTN08j1wlYbUjQEtnBDsPZs+VgaNlOxh5hz9PW6DE8+x0f5nv9U0jyLIHlyQ4xXC+SpZ
h4TG5w4wH0AMEbhk/FQ/5O9MKbIM1zlh75mMOEX7p1OBigfa59DgE6408jDv/VzJRlWTChuxMsfJ
HPicAqEX/ljfCAUlEzVhsR0J65biaFlUhWzvR2re7liH8YJzTfP+xqeI3qP3rRLSGKMJ5qU9V7UI
LxCt4FgFKJHucVnyq/jCTbbu/BMN5MdbEZZP8gOpaHWBtN2YVL2g7ypRhPqEnj3fqcw5B9BlwQWW
L8rDedMgR3r7Vv4M/4x6mLBNq4OcQnGMh2BDgECP1lSQHgpeqDO/OiWaBww5V5XD7RGlwzruv8Ol
i/AM2P9uoHR08OXClqv8508ntYT1GAr2bjf/hNTDri+JlqmUB0EhDLd8MXndlXclaitEa2JZ2lsq
+HM4A87smcAtjecMlfm6nXOt7wX55iL+sM2okxumcZ+W5vY0XFnfZemZyp5fxQLAGmzTqolpcYZB
eKE86tlbkEmGprF5uaXdM2BDSOpX6AgLnwLmEy3qWSUqwZtTjOEXX0HvTvyudDoKZhFzTQLXOaNU
BbDUzyjqPJoLYYw33+b+tuXzHcbfCKrR/HGU4l4TEYcdgsTpipRnWUhPcbdkcP0bB249KcWb2xWd
xRZh4biaOXqBn/FfNcmZVVac3y9TFFTnBBB9S70ZJr53soc7Cj6YkmU1k2fzTsv/jDCmd48cBzgS
VP7t/EONxUqK+06jcdOJBbp2f057aKMRu5eKYVvxWe5RwmtzZbyaxEhvrR7SNR5xzUTt964+nCn+
jGs4DMCAhb4KJQu2C+wzejP4o+H9O+Xhy0KExKNM2NYTYQQ8RFlzcVHkUrEm0nks9gIH0ljjNpnE
ZegWwbQC4mNedb0A6PXffpD7iljSbcgAfs6dcixK7450Xl1jkze60FvtnYa6+JdDWvrpw1N2fUU1
1EX5J2xvJPII0A5Whrprrkm+sI0PTIGEoFpZmPKLRABqQIxhRQUMznqUyGcJeFA3mW/LMrI1ESX9
fV+mjIGTN8mgAJPRf/CEmwEW+DGSK03P2IQxLm5IcLgSrHKw1bW9q8NFJMc0E/DkaZcLshYh4B/Q
jWHqPTfQHmHMLmJeA4U9cvyT1UhSeKT8K/q6Z/CRY1kFStGoi0uuoWuxJ9a0kdk5H0DY4I2WcQHr
GwyW/xRiZK6Yf2OTVTPByPu9OgpFSv8Nd7BexNxh9GwnX9q9OmgXh+zaO7Nb1GNLH9tXF9cDPogU
VpGlSXDqMnQNVvVPVRvB5MNAEOPy1kJD+IP/Q+/CUlZHGBssgjy+Q35L3hjQdW/JYihfSrDvHPIK
wcDk+LrMU4xsRMVahZq2TX/ylwxVEA5Dm5ysGsjrecN4+MVHZ8BaXzl98PyDAuolVskl2tCV1ukB
Uf0kXZjuvAPrzLJXA+mB7UpLm8f98mLNcINF+a2Gku3I4QabJp9EJUckcKvLeJMP5rxxTHUKduCm
U2Jg+dbaeMrXipqP89BH+8HsUoUckI1HMYa6Ejcli8VetFOfpcsTJBEz7BQntsYI4DnjN9W2Ntum
GZPCf9nil///J5nbwVUYrcV7lCIRHVvTYoyFhtAN0Npq34giGAtVisOPce5qjWOSPouRlR6ZBGp+
j94Noll4MyTzTLROqXkeo1JlxANxu/LJRCfqCZg3Sq8seg/AC2Imse489nd0ToN7W3c0XjVH4Y1v
c1/PwCE2HgIeSJ4oc6ZMKfdCOnDL1kQEEMAa2aarKbUY8vXaqU3FoLVGaY/MlCKVgqLeaW3xFEqT
OMXJL5M24z9b06aQWvAKfv30r33L/wY05dULTR6UiC4XgN38JJxqdKv5kxaga1Ln6wLIPE5Vmm6S
impMAV3aWotQWkGwZb0jdVOAp3TeKZmxdSG5pIW8YXpoGVvxEY1kPe9jWda4TC9ISKVsIK5McYK2
BbBWLNbWvwGz30HEeojhnTpeuVNc9Gvwv/53rtF+B+6CEcekwoXn1R82wN6ZLUdt1IZ4PGwmFdcC
gL6ODuWAVx8/Emi0unS7kvRsMhNt0xrc9HaWS+6riYm6ZgIkRHrW/fu35pWcIw36PHwVs/yrctqx
7N3six5xr4ZMG7Q3nGUNfaQKf8RpzRO4X0TLC4xb79p0bo/6gaUNGt2SNws5z2UVd3jyg/qDhZuU
t20w5BdiMNChBMBmpkus4QFfJtahuGwYKx56dyOM9ut+qgH+8PfoUMqMc5nDEc8TckQYcDr3TaIU
2kywFV1CILhVheWaVryQDmeMVXWB1pDDSceFvALxvrAlyMWOCK/H1kackuGLrSmMT/UYkAy5ATC8
/SnWcu3Tr/a+ffVcn7nPi99zq9oIITJIR1qC4Xzrtm28ORS7IC7cjH429azAktoq9EH/P9c0aRBs
wFekBNt1hsxbQ5TRlMqnjXvq54QapbxPmSQjph9Oe61I2hKESi8cF0/GRs/vEAw+aMUvaS2Ds36O
xVhQAOG2MYSxKyXrQTwUiI9j+9ah5eSwirvg3Z3DcVzqjWx0txd7H43OSK5LmvQFLqQK5JAJEFy4
LS/eGXbwwNc+WgcxZ4gRXS0q4tnESk5o+5Dkbnb4SBWMFh1GHVyQ+jBxwmWvwjptJJMS57SjWp+r
sk3iA1tPSHY0kZHPvbOznBbKeDD/S0ahKHaEyj4kqY1trHD66Yd6EoUv8vPY91MTnOuUsC0Rjon7
SUA+Vj6mwUvEm8Wx2qQ6ZY47+NRybn9zncuJ7YS5BsQIenQZNhCXJa2MBLVr96AqWyjwQNKE1q1B
ylM1tgao7wlIJW29fbQYBrUtMa0W7LdWOOAqQ3H5pVdBHxXh5j8UTGPzqKyNV+VpUo8tSiJ4XBpH
r0YFNHsK4xSw7lsz4kDbfEwy4A13PrjWmvm3Y8uSzDNVhjwvMLxadjo21stLnf6b04uNXjXyf7YV
9O0tRaKGzFC/Yl+72TKKIWd19532pcluMG9kkdv/n1B7DvQxsaN4HF1nDOS0i+Emeb0ePD5dqZX4
pPZdKV1cZAc7txxIF/nsL3hl6yc+m0eDEKTMhkPzqUO/ou2/5ZICQZeQCPzyy1sZA4F7a0uAcqtQ
M5j64ZcLTC3vVSRp4t8hepcmOF9ookgG1JUVmwmuNky/BxstIA0g3kXr8g7CdTbcjXP9Bu4Vfw0x
Gp1+3tkRRdGDCGCwwv4R5AbVFAamD4V9mX9Fmw6s1y6UEhKupB94YIrbasV8xBTLU022V44HZO2l
MLRZbcTk2UmCGjHdUhgVByQDODGmRVgzhNKcxYEoS1pW5dqNYo2EzIepSiiYQYpxfNGrKUtMkYVM
T5vi7lW5fPUN456ck0hv6NcQEdWIe7D0aZGqbHcqbYLKIGcaKWVZmsAUNdrwCLfHGItsIkTBzGkY
lKz86HiodDMs5heyN3MEzQbkKVzNhGV0gyRKgNNE5GqABx3WakVkbQKnhY8C1WOD3NOAua1be4+b
V7uLb1DUx5v7ZSRUlOBQMIZFkI3MdMWWYB2OouQKUwYNHTLDK5f5tCvplwTnRsophMZHKAaRafIR
jwSGcfNiB3Yiu6Z6VZbFPLkT6aNYVI1gQOamH/46tmru0UdIkkR/+RBjk+4XCzhGO5OuJNdD28N9
tddQ6W/29Quirz9I5OZpesS1UNz6Ki+ZAe/ROx6GZwAPiLFdIDvdqxsRM+dIl3/xw8GsLtwAeOaB
+t3T2eVb1k2maRr31BGrHK83Po7/PcHtpvT2ZkhrY7yL56Zauk5o3INSO94YZbqB/jcu/0tZEeDW
VDzHOhNOwnBbIAbc+6+VL/RHo4mwAbV5hM8WNtvULVPekbsRlDgT3cCGSbM9rWwxPmqhm+mMH4ma
+GqjstIE6Chr0V9r9KzOR0F1ZKWLWeAmnafB6l2+tfH0xdNjaWCQCWRYgujsckNiy2v1Rvp9ZsVI
e7kD0yXSPi5Hwewxl+/H4Nb5zhGFQr45b+DOjRkeI6O83HoQsgfM711GIs3rBdNPTPoCzW0EsBz7
BKDVvyFkd7hxvmbTQ755vWF2ZQfqX6u9YDAXHG7/aDraUJtkj2GYuxPMcSKa/vA6UrSvgZggiyn7
fg5aMYvXs/fEXa4iU1LHfzhKLvDf8pysHPwE7eOyvHghvLRvtlXBmRd8sj8Trr/haGcAKlenBDMg
zgj0FOEd/9Fy6DrFVXuY/2vQNj+Q3g/G05huIPfG+IlFKsqTIk0C62eJno+EbOKJJcE9IFdZBShP
OB1pn8r1W8S+ZDSibcFUnM2XxbCXH++3FsjEbrsPpyIOTZq4uLI/p8lQ/VsoMQdnR/QWyGf/L7Kx
ZJlfOyOtTOLJbxM1HOphTGeVlD0QqisMJM9tkVSC3oCFZAy4qI8rn3mtHM+45w5vD5GWz+iKvQ39
MGHMdK9dqYdjUv24XFlN/9QqZyCszs+rvKctMIC7d3anR2Q7Po0h3JwQd70wXPZIY2TkHkhbL85T
Y0/7zLTryvL1na/D18rp/rTyqXi0z0BHEn5qXi/Av5DCLkl1g3if7HfaboJNRFbrbXJbY/o/6+zm
zJdZeK7cAjCxHJHwymYCcSH8PSffkg8pb/tW2BDRHcY8cPEMmUpmA0ZZx15gNvQWDLGJ7j/t3p8l
vucrqbT/vdLacFrAmREqQSr/VNV+sgdLWlPj3W9KuChGoCG6rNVMxZxdQxJJoou8/u9pLxnDUzcj
zLSnSrMgmWiaRLZQvesHNKvbmQ4dNZJRV7+0RaxJnsUQiy4jSVTDrQZxY3eRlvFsiuVIwN0IsNSs
mIORCFm5DBGxlj+C9s3Gn/DvlctzUnUtzWDTs6UcRCU9+bbDJ8ayiem3161kfYo4TaFBsvD88oF4
CtRFtwCeWr5LiUYUZjDUr09d3g+Ab/w4IvvMU6pJxcGuQ4JdCGCR2qCydtas2/1l/jbGWzZBS9Qh
44frE+jjLUVpnm6Z87f6Dhy+ItccCxIEfI7wex6sTBeLPz6pYhmBhYMQSIecJkOVITJJm1rU5Rc1
SlmbprfPh5PxKeUJNGHL+nGv5/opwbLrMztl1qSRGVvhljvQ9N/2MKLIvJ6rAYKLgp0Druhadvax
mAgqYo3uavsvTTGLIiLcLpwGO+xnL7iEU3jub+ErPSc50lxf9/VRR1F0iqWqbR/4ESs0RCN/cNal
JTYejjhrVyLgnMknzM2jz44gW4FaAavJx9XYh0GtLEhjG36f7zJ0KBMYVThvS/WfSLUXlb41Sxez
WpNL2Xgn949ULhUTbuNSaYcWppHs5RlZ1ErGgZisqMjzhvS7iXhCn1DfJT4i3+m9RxzvwhmdNh8Z
STbCGMw7coCEq3XM/9e2nhfGm2oPrn8z7aPTvXiQjJ8Bsq4vFVoFU9yZV54ySWRvNtRbEI0jQUgy
XDYwvikoQogtSpc680bVEZqBvI15ruD7YwrO7wURcAMSO9vNVPcXe1y/JpGP9iCXsOL4KXU6G5n6
khr/R9xpNyEem8hm7h9iyH3TzdsK0V5wGHotDtMF8YvZfpNln647m7krk6O8hKEDSjxGEAJljXIa
vBZIj3frimGN65OT89YG2iYMmjSecXTP1VFy7yWPfW9ZgHK9z6c7mwsr8r9jbBjstwnk7+pEoHhX
et2KmxVj7Ab2FnQROgCK8mJn9hD7MKOXwyqF1u9cJHpr47zXbTIKmwqC2N1gC9VzblxZE+na9A4q
GyEhdrd2ZozbNIUZH+4cwr97UR97q807lKVlHpVAzdnGGHnt7ntwxVb8TtrhvcdtrzLMwBDb8LfV
bdsnsgLM9aVvYVme+yFT31/O7CG5eztf4oQ4z9coi4sWmXUY1r/qrSo6zfb9vOOCOtKsgBoM9o+1
PBwKadZjuNzXrYuALcuw3mrIOp0QHCfkFwz3ZhpY9N+pPJhtZQPKXE2THSiDZKwopvd1iLKwZas7
FOU8i/ZRMkHSjuFd58UL+xoFvsHwpZflI78bs9T023uoNp+USndSrS3x/zdMs4mVDVPCTF0eCvzv
y5zzoKXHfDwO4sMsAsJcjqPAVfAPfResByQvy00+n2S/QuhswCGFKesEkmp2PeXPvpLnvplIA6QL
GSJ3G/ugtbZDPql/v0qBMGyKPZssWokl+QwhwWeRTm4/HAXVHuX6VydpP8ASAtQ8FNWCrtLq7Z9N
IkF5zu+c6g+LRe9mcSzbqJZcTTA/mVjWGN8c9bdHVFpBwbKrfXTE1bRgsGJuz5jXq4+KFd1GTiv8
NayC6LglIjjD1TTBcKOGQT1APuYtVrYcLhviq8zC0ms0IfT3K6Wyq1uZa4TL2oBqJbBtrHrTEU3g
zJNXbU6cCJ9ElIAB5OPOJSfkcMFfkTDXyixf/yyY/Q+BIm2mcRhofY/TsxvYT3sEo0Y5nOo/cui/
NH6cQZ9yrrXPdXHZhMRDNJC/6LX3nAvai/gTrzlFDdusZhMXz9JdHf/aSouU991bF+/OyrW0Ilz1
lkKQhYnlx3Tn2bx5PbzVO0g3uG1C8fWDptcXtwcGOHbfb6qOJ/wWkOvzpW8e1jvbRqT3DBpGNtZl
aU2Aev6WU4kkk9jQL4ED0HzBWJxFglnmNYix54/QsUiGHDT8VrDvGix2pkazdJJGABikFXxOXOfD
wn6wckWPJKhtkge62RB9Hq1gghvMzsHcpYdaFzfnNOehdb2hFQK6AVH6cfaJeqt5szLvGC8lrmv4
L1Om5KaeF99dQDL8w8donBePi7Y1gxrSsZQDTTBqS7LXrt75zE+FBh+tS8LLF2qhkJukYmpde7V4
W5s8FgScmKE+mrRNzlMHvXXQMG5VKNNmoGkd2KmjkaP1QCgjjECUz/j6/1Xo0zpFQTSREOQLuRIc
N3YbiSAK7xDYkYrYrZBjoTxMMFohVciVl3un8REoie/xPWRkoT6qGlu9rlFNUYaoMSCu7jtFeYll
vpDV2Z6ZA2fuOP6KNtrtiOGV+LG5AbOct52EfZGiumjIKMOUXRt39iKwEXOdVxtCJ/8FR3TrDxD/
uGoo0NoWG9qrtxqUBwhOikUKM+LLU8LA2cnsdhOBW/C53L1LsSBW6JROigs5mQ5whM/N32SooWiC
RUmyPTyIizrwJCPZqLDP+duq4u+cS0reSN5bK2z7RW+BJ+rXlEaB1Tpz/zMsuln1lJGvsJ+HZEGg
dGaEq2EPQ19/WfZh+MNxsRakqGt8T/BHZnV/nnf+TjjthWzemr/ko40sYsnrxYXH70SXYyQeaQ63
020xzA+O3hfRs8Sgf8E6uSwaZqP+9bXciiCbyUl4B87dMcdvDAdVMc6f7CeUF64hx+v45hJYFjJ8
jRG1jo24QE/Dx9PUWGqRDsiwMjgKp0R9Zf4wBXGZg2LD3oPdcOVcREjWRE/xbVINrD5Si8uCM2Vg
ZE/vv3ouegZqia9J++KYmoT65qrkE8ARvqUZH/LdI+Rs2S960r2gjij+oST0DDqa93ye2kw6Im5o
bU+2BBA9fzsHwP7BdagMA32TGOCVf+lrF2VtMqckkg1g3e0Joz5vwE1u63zt7jYSshn5bTA22Mss
cGlR3Bt8HWbx2VL9TMxa40mrhBpS/yQYeZaLXim+yqZPe0NthvNglmuv2vP2f8vG8fheaK/eCNR0
NOazBVfDlGYmQCaq2YrOrAxtJMCp0/FlVoFxHXdmFxDIVukdT03lNJa1Do2+G5176mtSNcB/hEuc
TiQr1IMyY77ergD3MqLw+NldyKQucygtxoiGtfwElkc/bq0NcIpfgYRIn5SYouonx9cZQtcF2TTt
SdNodKG/IjCdI9Fr1bqRiSqFlCYNWxgcePhRV+ZtalqmA6K/DnKaT8I18GVdliwKtx4k9fw8s2FA
6+FpNMLNQSYxhuAghmjMr3lSyWeW1tGk1hqPbPprcE2XLMB2J6Zuva2bU6KwcxfSvCrYGDfZ6m3n
4I5p33EKJ11zV48xAVl+g8uqCJy22mLX+V57cDRMeDHEcW9Aw/SIHli/yEm3YNdt50ORchLTlNxC
O9ElKVYDvyNbJmE6IUvg7dn6PnvSwzAbMtA9Gr+47Ec70VAVgW4viyLN5DuLypIWdapAHfOteaAE
k1hmftMqNfwp1kXlGL94SoGm/Kp4G65BSAgwzxpRs+kLwG/5OiS3wmdbxt9orLO5QdWd3NCDAI5K
8++grAtvjGuZGtyjBr2le2wX3WtyhwKBOo0iAQOAamYBdLDP+YEIa/q5G33ovswoGwEra8gupnW8
xkpUEdld6pl4YTF5Je5Yqt7KuEJKUjYt+zQ+NDuA1/4ZyqXmIOlmDgXCSoU8LvGCB0q70Hlsdq0N
Yr71RuB/q6IwTKhnYqQUFBxlYvdRrDCzCRy7QK10tZQtqLvPWbTLuwQ7AHU/V4PjJy5y1wnZ3GYw
Abvxr+lkZOpzLSldtX+3eeXDkrMMZ7189SfQbuom3eiIn0aq8tD6zStQnUkgxLRrBpB0SGnFLImw
U4RE12FncNBB4WwAxhKDbT3EXG3rGTxXlYn3Rf5CSst6W48XkF6659c4gK4fyjyNU8gIHHMbKuN0
Y40mdNLWSIV0oEmmpi4Dex2pzqcEAFMZuYm4mo94v2Kcsyubq9dIeD66OqW7ncR+W92Vpx1szBUE
KFnUvEuBl5oQcOF6Nb9guh5zusV8v0j/qelUGbcmS3ZVRnzFDG730kNSRdiOdXle6TB9T7YykObH
wHhVbDZ1G4gqA9icIj41oCE9Rx3sXFYd0TIzRNSW6d7OIYiWG/wODrVV7+O0KuUQw1BBrmG5z05o
6qlM36+B61d6rEhT9KTmvrxNap2EYDfy79CXEW2/MGKp5c9jwPhos3WpXIItkI6kZuawQlyJzTee
tuosn7mz756zcx5ZRLS99MVCc5bREQlEFJYXIKvRUrr/BWrb2lpHDKk7b4yipq4ldmoiyZnSRwSq
7Yn7eCaBOH+aeiGjhv24O2RAapN/fyJ2IM3r6buSQAI4WMqXQy8el2mNrirlcBfxJTTpreeaNTRM
FA2bVMFBnoT3/X066Ls0blflgjTaGCKUEhu+jOYEb1o0pg8tXJuMgLdwfpt24fQ/9sAimbJIxIhk
Ocp9JVemEwqS1G+knyfbb6sh8cDgd6j9MwJH5G/YL4LoSgllvAjlA4orRzK7mkOU0wsL9iaF1pJc
OYzxvxFLJgpbfLNzckM3nyhcbQ4ZDYPf37Zo5djFqtPDnHXa0Wt/To3r0IdruNQwO+Kf86mT8l6g
w1fBsLJW4xIkdhM6X2XH3ZIFqEEp5CR9Ol91a9xBEHs9+Q8QRTEjNVKR6RNIw+O6/uxa0t36CTkA
dlYrl605+t9t98JkIQmCml8/dj+AimKwGsWEmg0JVLIy3zIwdBXzzeR3TkKLiAINnfJNxIou0aCZ
IUbnQ5efOoznDjN/HY5k1LDaSs7mwGxwx5XQQ2bWNchpQcz+I4YhltB42afm9/RLs9bXGTkzLS4i
UXjO/YduXLkZWQKBUutgsXGoRo5ORkhHciiUow51Oz+Twj+dsZah+3pKQKWzYFc8G4WkPH2/rZv+
Ry4B6DKh8bT5BnEcAiqkKV0ehMUZarqrdsAME51DVstraKaZfMxMyHqLucT3cu3SfZ5vbZx80smc
v99zzAxmu1rU13qhWSlnTWFvBETZiLyXWBjsbnG1oE1tS6uPJhxYhxw6tix6a1AP4i8/ATxlDRvl
pYVqhDIttW1uol4B0lfLAoPZJ85Cbgnj5BfQdyQBnSKhLg5b/fo3xDwm2ViiNetyNJxvfcO9CxFL
39/An8jO7c3gyJcE47vMbZy4adHYvMv+Ysp2pQ9QqurVMJu5+cZTBAO/VEcTejNhAbNAEUibZ13/
jCWB5II/6nKw1ejVLXdHTGpB84xtShGstiGyApeRiS4plGnJprLNoXZBEURiPvSNOR5YrwKHXezK
ijjPdgg9t/m1+MGlFztTusAfu8CD9pApDLgHEjZlIk/1QveVlFTQPEnimAAXr30nW7ZmvyV/1tmH
a+8SwLIslYQrg2WXhtK4rU8ns1QYxTl8ms+nf1Ys0TurxSWzSgHX18GW7R5osLhbRluN0S8IgmZM
rVhsAxbR9vmumCY99IiyuuI81sAVSp0S09FqcpT5Q1BUNj1c/DUYPgKMlX2n8GaPGMhlF+cGWaEl
uU12OUes8nbYFw28GtPULc3KI/waWHGL45srqvhg497svCWw8z7QEq8ElJAemux8PGGqTnsaIGtj
+eQ2aTEGOO5KV55ZCchbSAflvpWvx4ymEbbQQ8skXvAlys/YhK2SpVNC1NmvFL8Xe3VGdXbO5kw0
UGyGUiv5mln4eYWfmBnXLmyzaDHtX0lm+qJfIV2fUA1RPWUZpa0V5zZShGA3e6Wj7AMYuAP405Et
Rp4jVcbLwdalK3JaA6kDeNp2koh7G3Yy1nPpAyrG8+ha3tZWwixR7dKVh8gnKgaBJ3meLwMjtDi8
bJQs9xCvQCftgOS7XZ015R1Fvcpap49tkrVqxya98TrQFzohOeOQhlkLOfisgDfVjnLL1tGWgL/L
pLQuJJrWR0yLY/RXG9/CwNKCykK/LnupnFgmzv+RawHfaSsgXqDuvGsm5RbqF8H70PsktQq/Bp3n
526o4VTI/7noxwb1ku0W3DksepOopwlcHP0phAjmxbfaotBAWFIBpSeYtMKeyPzV6zquKt6CKl2W
/TFgk+VhqcN72UJ/8xaaMXFalkwSKh0V1GouLMlwRCDTYqwi9HYS2bWTNF9pSt81zfuFMYvyQyQ7
ox+t5zPU2dYwp3Mla3JEEk6scmFiebTHTHFAN//c1+d9KUVtNUjRV+uFj2irKCmxe8KU86nk2q6V
wQpEt/Aux89f0vKp1LxwbFQYNQCXU/KcxKPge8fE+9UdcfUd69oQTIKK3oAoYc7zzP4F0xghzLKf
OwTI4dB/7LOJ2PbyWg5/GYjnpArXdiO3o3ibQPxBXF7D/fBIh/YvBMOQSQbUMA4Rg598jRWFkxag
zJIrs4FIvORvgv/5qc0C/KZpIb+kcFvRB7Ikusq5Xu6GfG4ItVoSAjd2Y6f6+vkmQMdynnq3OLEv
bYBUss1efahwnFKkcSofNKvyH+v3xzeM1RTPL8jfV6ZQ/CUS80SuTlWg6N9+GtcWBws3KqeQODNH
xsCQBTPvQfO1WjhjIuy5MFMq9xnoqiRFMIEiJUjcTt4Y+r0HOU9/a50f87ZGP+gPuabcEtpzE51I
lkgbJrE6T0DfVYVdd3wJUSUS11A+vdf+JJygzGqVGAKzf9qDczl2J2HdbLcHN4UZMMTdbY8RcHaW
KSXwMTtNZWvHRs6FnRc9nyOxiIwMcLoOpIG6taQuOHT20fhTDH6MK9lT9SVHzh+LjSKFY9V+ScQJ
vAIxk+xHUi3FzIIfADW+4uKWb1m/Enm8s1/03sxJ3QXjAh8UYDuVeOJjId8+sbSGqxBk/n3mb5PD
+qcy/GTg7CBXT+KE6BwQsweqGBc6nncVElXKObUBAEvhVITObgyGQcDhKUK0LoL2hFNMxwhDN4/W
JD4sOOm+1Md1fPqmB0KacgNjCGSOazhH/OtpH1qKY9lUqEnJXGVhXRVtZUzfcE80VW9x5dYBFT96
7K5ZJrH34knvz5qSrU9i0pC+UHu93ggRvkW7A2ALlfmfva8nSIK+qTjgTGPd+EvD29xMWbluWCQd
HG8n5H1x6njOxk5uRh2Q6hqje+eybFZd35E7YOL8jT0scdpAGs29GyowcEKn7Vpxz0aH3hlS0Fr0
QGAvMTVwsJMi+h068sc2icCrxj58BPXNgF18GG5YR4X3Bb4ixAwjxp4/qypSsPts1x8EBvrY1hw2
SngiZiMibsQxrn6KlF7DqlR1t6PbECpJpyD/VZw/J0ONWobiR7aGzM2UrkCXozvF3jCyTxhnsT3m
Nb2YQ9oI8SlJo9E82ECdlfgSR7aQhPXtz3dUJ4mO1ydCu5n8VafsvTlPhw9JihYK+ImVB+LTlQeR
YxeQpsNbmq15yuOazhe27KDME+NzsInQPzlRNedTkHDfccKEfh8/jKD17/aGNy4xujP5CM7ynUfi
rEGLWj8HRNha0c6Eq1XbElklJqMnA+Vsc80oSy6mLdisggYhgJSi3Xdg6JVUhJHAZsT9eq4elOaI
PSYuTrZdqxROGLfuKzBEwHkFLFVtbz6+noiJsPoQ/zc7ZYWguVmgtlQ2xJxwRazT1VXNMkQr+gBX
hH+sYr8O7Fzt2sRwoHomj9TNbF/RPS4X32AE63JeJGP3PmHDxkOq9EOOkm/dsxz33LQ7+Ie5ji9c
DkJ78jKI5otpL1puS7fHzOoHo7+fi2gt34jOIo+lcUeToGJDJagmltgO37yZBcmY4RwC/KBrqJBa
qw3hnDXQti92GCTnIJXywNwG3oYCJHjKNSt2s6M+qXlYaZ6qpO9V1wrnyCimRngb1/GXIn78bj/R
poT2QpQ3wP2QhCOEhYQ4cFR4efSzeovEWblsoMBRQ2uIY104KATN2XlDPdsfdjBRPD50FPM9eONb
JHgO8Ix1SZTKtKJKcZEipHPeeGk0HRo/Teiu9HPvP8rtIyl6+hQOwev7OCswmuKizs4Qftm+zkiw
l8A0ByyZ3zPMh40+ehSPesJLot1+Pb2DhOnvYYSLKp6kKbAmf8hyGc/e2MITdGZxrrF8ep/uXKBK
RcD4M/HK8SwtK2G5j7OUHsoBsNEKRo8lC2DUWZR0tpI00A6aW29Q32HA+MUnwYnV3gAL8qb/2Aa3
/ojAILhfAOqqKA2/0zp78r0vnezhmmTDms5rVfTGEf13a753KiiMf9Aqx5No3BS7squSwgIJLAHy
bmoxvdKOwaeFjan4gX1NZkNdSBbO/ehzqgOo3tjhPju0iWaK1MD/vuvnPt0qNAjT3ZHatybNY/Lq
VtAWYIxf0M9VYEDGo947yEV7yKFPeHwZr1g64GUJpuBJ/V4uG/xEXv4SQllUuC7ytvEHvlkNpZbw
NUJ1dIqplisqEBddkDc/MNFmqKR1qoa1zc2XJUSuGANqKswGZ1noqNDLl+e+aURegyfXBVvJJmo0
ki8uNXoNorYdDwj1rdNdqOoYNsbFTYzlGylwdG9eAKZL0xeFx9cdC3j77z84HURj2WxZu0OJ/OqQ
BwyQVjrIV5eSWilc5isGKXUkaM/2qty+AkwvQXTWeYeiph3zPkOeWIgEsKwxM6IXmBArUU3qeb85
zGnDtfHfcrVbrcsDNzaDtbYWzd1KBk3XRzx6wSunp4dmtJQ1bTnmIHpsFfY5T44bkyV65B8jL/f2
bRPbo5rR4IBKFg/9z99f1RDtuk1M8czzaDpJzjYhG0/fSwicq9HagVtvsu/OZ2fWha7NlIvVc12t
MK3Y58q15jaf5j1s3cHn7PthFFgZiTwHij4Ljz7YoM/Ml2I8sox3mNznxGrTvkgU81VbaMO64Hlm
QzddEn+C69tChS34ssQeUe8hXTjiQsQcZyolGA+vk4gBiH0qE92EmYFUopRXF/USvdlcI1a8ctUS
3BP4OoNd6xlZU9+SiN5RpvgMC8rOcg/Xwz/dhgxiLu4NR+2WdQaQG6DzMW4vd/NUXOglgBKXp9Ek
nTJifEuj4s+7I9F5hgEhVanJFN8V6g2mex4dU4NLm+NdqopS98/Zo/MA3wULTWLzC8/qUkkeDlwz
OdsTbEBPAH87bH4uHL4KbkS3VnUBg/2Dlgj0CvA4/dqXIN9HxVQ1mmI242vVStLGZALXywED5TmE
JqxVdk0u0wqxXjje4ydjvame6o+y1PYqueLsz4XCAuVR8AEAJitMI8ntuKA/U33mWZooJvCi11Bx
qJsWkscrMUjF+epg6s5oooUO00SRufkWYh0CtqrCvp8dOpZdavfcWVg/EXNdufWwxP4ttYVWtJFS
IWoD/M8drA1ixyp3v5pQemNRIqPx0Mp5ylvWxexoh+jhlx1GTE0jD3PBEyZPibOm70QuYV6TcNdB
m4KFRNZj7kkhLMOKcl5u+tGv9N8QR9V9GUGceIgDAsz+MTOkg4/rGpboEHG3rHYo7kYg1HKBILMC
ZqTeNR1WXnlzDlFOs5zv2GMKdrQKsr/C2QHp8G0vOwasJ2KzDDiSu3MskWpMmTQM+GvUe8vowlV3
n2R3SF3osgVrs1JCo6lMfuMmUAiMGvfgKXKIJzD5aFEBMrFJhLZwbAFH9cYQzHqP0QN+LJmFowKn
EYJg3QpQlzi+fA+7g6z7n6P3IYsUyLESkMcTWcUCd2fx6LpUBv8/BL5qsc41V2D0E8j3LjREb+Pm
j0KZ4DG6PTqwFyBHOFceMV7yWHs5D0p+KRguLfJMFTWZChxOcMIjvTYesFJ2HKIOpkg4/npvqzNQ
JsT1dQc5AgzXFb1QQb+hcWLMYsLTTTuekcyIap/23wjWVm7fwvstK15TEzhxjJSrNqfifo3qkwAM
mgC/CDPErbitR9VZi7WsVfboXH9EZzfG+3hHf5Eg0lNf1m/oamxJ1/aMXO4HyB8743bZu7RPV7sp
a0Sp5QqrzLljAoYqeLdf2h8v5GLnBG+RhHc5WvvSncqPaNvzwqD+CHuqsyocSnDtg2X0ofiAK0r+
Q/tCZgJ8t5FozAO1p5v3PKXxX/r2pVyH2rwhq7GbTbz54TIHqtfdrbSDOhPvCWbjcL5YXdHM/UDm
8Zcgdhb2A43k2kmlvFdf1l/ddObKZEOpOEckxDTq4uhYnDNv4bmPIMdlEjM7RmzEy5rw2+nIkWb5
oYKf/wNc0Wsdu7Kv4FfvkxOfdZYyJtxrmdwtX4vcsFaZVGI2dwn+g+6unSBpRsHVMgF/GcFRaeaD
Cihj9SfGQ7tWF3SchFKHtM9B9/GP7oE0e1MB9YKR6gwSMiTfypbjgpD74lMPaP7E9XU3u+mLsfiW
XJgcsNz8hcq8PuxGuqF397yVd9+xkZcQD5zex4Qc8I5d0S9tY3I7FNnhp0ZsD0chPYFFNc2qXK+P
nNrFQahwFO2/wwMV7lmOxFRjTR1QSx7NYXPUEzAwwkKFkN4/nQez0APwGwEblZQxJ87pQiWBnq47
tQaaVDWdcRPlrBW8tFbDF/YR/CbvyC7C/SATJW0O4Htc536xlHLsqdbrdU330UA6nevh/R81t2l8
9Mo7+jfeY9jeNacXogVsVzV2UNmAHScLzfJa0xlnkty3h/DvQG3Cp/4ZpIecKZRPGYv2g2LIf78B
3SmSP6+lk8vf3c3kTJdaYb/+4jBjD7t+sahAHgZZO8rfuLKLCdmtUZDtVqCYAnyhbaIvs8E21b5K
6MQBrWG3WmGnAe8IgoaHbq7msfKd4hezDfIrCUT/YDelOTBTL0ffdxhu+VUsNOwHHvucs0Nw3Jrs
D3u7lNB9cnBTa5DJNRFJ0TeT280Xn+bwqImPyHcePArAyx6qpqIxoFWnk3djc7RnS1pJW2eLTpuq
qJ79YI02C1jKDgOTtkT1LTfk/UnYLuJBiGpUTOoAeA1TMNC15YT1N5H6NJl0XNZxY0YkcWFRTgJP
zIw9bhw5itxfmK+dZ2a1qGLdmHjY137kEX8ih01CtAQzJ73RPDpHXfsD6oZfgKXXTjFJXZseLgpO
nS+mWaAsULmdfDiIeJ8oGhTjyE/P84X7lCL6HWGIzwEFLj02H4bghN5SX+qm2MCUkY4ta9i8Vs1P
ON9Q3Pl0yjO5eTau2oiwOl+gJMvtbLSxI4/bxwMkT0DZ4Ba7ilGLe9C7nTx8QBfyq0LmQuPMnApm
133fZ3rsFfUqEj8FwqsAvDBldzx79Hlj1vNskGD0XSVl0YepWCrEHDIaJmL2G8zo1+YtzVTkzCAs
1YlQPk1XNABdFjt2dGrbmkkUbP2VbFZtpw5S8uvQBowc4U7mrMKoiqL7TB/XtY2XX5sIwaG1YhA5
MBv/XClmIcEyd7CyWOVA5ze47gDko2JagJo8s0cHlitrJWrhdXDxHPBsb1IteoSTUVedqD1uwUez
rlPjDslEvvZySzoEw9l3r9I/OWiw1R+XfCGQXi5xLwNyqe2IdCvwaIq2cHKZBv229u6qFPFpBauB
O+iRKRS73L1m77/f0eAVw/N775F+d3Rjy+3C6P29IxFxRZDWwx70GvV3TJRUy7WwRSJQ+nNKeeTA
lyQownPuWETBezv02x7L49HdwKOjqEXAV48Z7EPm0Syf0pEl8qJhgbYTk9tVUgYxkYc88ZIO9IhC
nhL5+traHiRLKkT7cGpdk4E1mpZU+DdtV4o+kLMzlTxqCM5MmorLTXVVp4fhOOlJbN318v6bhOTe
BeS2V9ufAlwTWrkOCeNRSXI4w2Hn2D4UcOYgocODYzB5KTT7fXsLEzUBiqRymno6XLdZD721bb47
rqzOAffouicSTkmCJL5aBTzV8zkCfHWugFX2liK5K+nCUNcu1c7kB5zj/I7yYaM2j9APBXd/MB4U
s0QtM0gQUa+vGDmKnxEUxRGDuQjx8lElLZN37P2q+mzR8+1rotqsX7l9gE0MY4fFmWcifzZiK/+o
foqlaN5USiImp2PWsfyWhv9WkSMNN5eUOpXkuT1rK++rbF0+90QWpkxORss9YM2ZGNg0XlyH6XpX
LRIMr1405T5ixjOImQqmTZSHrgKu65ycnfoB7MqkwgktoK5/nN4qN3djEkO5X2hi8r9GUedgENza
Txm04i/G6LJGqQMRgmqOvUSKdupnk6eyzcwgF2eQELyInUWywCNVA31DHiS8ChZFZqIQV3SOR+Sp
FW3xVEqZmV60RbOqDgWTn5RJ649b/J0oefhF1UWZvAqyda9nkHcP4CvBA1KwThN7WjbG2Ja0AJ2E
uyw8hiwjPL+bgEIAcbnJqSIy1dXKpbLPxxaWSDMoBZ3seeX2S+OtmxbHbGfUpLMNG7KsliCodfiW
PbQ0HzPWHboXrFHrMUxQQGnb7QHBQdd5rZDPGGVa6AMkFr+wO6e7aShxuNygFMCGpsNcdwE4n67D
/V+sSylYXugTOECZfnwTXi3ElZgBjoeK09fSNleKt/Ys8vy6w3pWdYI6v+BubPlMwd5kf9iHrwSw
OzxObLfhmQxso9oP5h2eK0qYN6mwqaUeVuwkTQ0PG5IKruYn1+EX0szaxBGirMYhGsj0qpMZM4pm
Ojcwi3T1tuJbiwdKBbhzs6DbI/5A4ragY+j5riDJeor7AhjCiik2kJ1U21VkASscAI8APt0rt3kW
vNSGejF2mYlUlLimNYTIeboxDTIaS+ZaBiUQUaEx3dwDDydxXhzzrG81uYPBYTHaq4nIftyV2Fse
4F2aEduh6u0wGjmrIHKkyzANa4KZNiabTqx8fdQh7dEIKuumk2yuomoGzD/NmyL4Uzr5iQ04Bmw6
g5pM+M9EhGEpSDyY2WyvcGUFCK4joG9Os8gbdw2tbQ/+DqYtbD7VFi6pRxcwCy48h6/X1bFWECAx
vw6cSKe9vyms43rwjj+i+2B+95pH+7ZNmcwi82kZQDQe7Plp6S3MNfa3/sQs8C9BZvPMpa4vlgI3
d0DBu/APLHr7vBDaNLnvmF2oF3ZkPqYMSiNIeaKjR7cha73jxs+BbQjzSMJ9lRoNbd9fvVWUXnug
ZSIDqHzZddFN04btxYOXVkZ2JUk5mz/9H2+dsgU9Svvpm9+XMhPIGW0SWbDyIgkbMtmLxwrN6MyO
h042jhDMzFOA5z/nF58GOJFG84yKv1N2xBDVpCN+EBH0NA0o6ovxyJjXtSey5MZ65RUCPPwCVW1T
A8O7dyUdwZDbEl7+KAzy22hnrgv96nOj/JiJQi2xj1QbhDV5uyJMBTtXv0XPtuQUuX2klTPqfcLH
moI8BC5gJBxqBvyiB6UrNKE33hPtSwXDLKbta4maFzvcuNjAqjyHV6119tt/hJ+AzZNsn3itrWrS
uMN8tUCf1oAxm+6GRvyF3giA4MhYVIcwvnFTwIss1WbkZvYZxEyl/r2cAJ8NJstdEIRSliCN6j6M
3Uh8E+K7fCeg1FrVlFcwtW2tA/YibHtX2g1e6Hq87GEfc4b6jq4PbVKkqkZTZCMmOPlVJCHUuFuO
Uh8QVNVP+mgoCtOu0vyXsAH9l97flrNpiF0SkGphl2xP7zotNjPlonKa6ZejFiUwnvtjLISop1mT
CJznu7vfjiFNeC/XyWpL2M0W9jYECnurbbnl90PMS/jOvEoCuMks/z+A3WaZzywSCg78OLuqc339
xcNYrO0GciLQquj0ZVTQdmlt/3FkAaxGs+VZdfyitYjmv5azmHkHrMOoqGmUgSp82DrIJ3tVwF1m
lfWRCZ8HdJEK3GTcl0Gwm3PSgcNYDlPR8fN9HEuAfDBg6lurg6i2rgEmHhqRb3XXAe/LCJWrxrDb
PhEjKXneTwD2eBiHRqTUK7pZwrhM6XpfB9xaIHsdNJ78YlwWi+uINX2Ei5j0gNqQWLnpwifMzR7k
jCb78I6RLOcq91wIjWqbUxCMGsmeDrpy/g7VXkblshAytcKwa9APwps1Ng7hd+EXSo8aThK+qUfv
Acafq3OWtNiXS5NFIv8jjdwireLJ4ilLJXCw/w7ym1+LB0WeyhVm2t0idySvBdnOKGNKmHmPfeV4
PiHuTC13r7GK0HgCbZQObMZyB6YlWN1vxPVw9HDFsqJKP/lTrifYrHQsKSEEFPZQFzzBDdUCObgU
DWQN3VkJxkJ6135qx3m3OrD47fUIW4l8ilmWGJqHVoc4PdhW4SUkAMQTtX9KiVp8Z5gqpKcDorqu
8ErAg8hdwQjctrMHtMybsqPrjGffvtjXvVwuwdZunZMkKeVNLlQ2xucGQRMjOZYcPqzl9Tw3lFCr
z5gewX4tI4ST6EWfsHmZMrrQzAOYQfTvEKhYt+1WAQkcQTNkWWmsb+ktSmFY233Bb/hYQ5iwTg8Z
OJACVe3tohDarpoggIkWC8l7MXFyPn2nzEWOi7LGkkrpDXPZgnh9RcV6MUNH6rxTywrzk5PyeYBI
PBsJJkEv6m2FrE3fOTP22gGrAiu1qHoL4E6khw0YZUOBlSZYGv2W2guGKFv5k/XramVN/rApkzHt
B8ICHBygo1ttuj6f1L6WcGopXNGsHwYaCY6RID71wLLQlOHzGj8ODSEcL5Krym3Nx/8Wz2wjPlOz
oGULUj+GkvhXBGSubNUeFC6NmpZgtjLjNBtMWaAbm8npCGbFSRjnMUcKM42ljiuK0aw0gihnf6/L
2ZFBs8U2PfM242MBzPGbumgOT7fUGaaS3xVN2nBPliTysQNsgaVmpeTv5EZpraAkAXvTq+3pBYD3
ciDfhcAY4cpChR/9lRZxYyHGZRlc2B/Y9fvNdoEc7UMFTB4A87Zg7s+4blS+z/XiQ0uY8OQim/2w
W4SVV/iGJnPUYAxUK4rZsXcRAyNH/mjGQidgvTAEpcjWzl5DF/XP5ZVEjG00NqBDBYig4HYDpx0P
MuDD3gwH0mKNBK8MXK48F0/MJFGJnzoGMA89jLI+8RgpVjfEjKoYZCtpMVEm9S3VDGeN4JUJvEcH
s8mH6nYOGh2zpYuHS2VWwat/tUK47Gws35kH119WEm0SlJCO4QvNR6iEo/Q+GbyZKxyJH4JTOnrD
ZVM7cDGdWn/3deVUVp5xniCBMabBOi9/0yhJRSfbmBnuo58NtALXeH+M5SnFQqDo2hbJr1xpdFX4
9OstCXyCLIohsQS9KqfUaSb/jjXTwBHvKsEz385j7h6SFsvY2FX2xKU+LD4mzaoO1NHILYe26CI6
vyIICWzELjHvPpqo1KQmVZRP5v1xWY9x++Ar8+RmBuNjl4QRh5IN2DsqWyu76bflQj40WnutVJLd
0ysvqOYIKzP+wyM31u70nU3l5yhtM0S1gWk0aXAEWJd1fBn3QXimLOnXddsrdP1SrmRdKFQJFZog
bt4oMAX//vtNulLQcM9lgnO6Bk1pPKC6sGgd9c9gvB/AXl0s8VeOI4qZY9pFcu6LKvFLOEL4TvHM
Me3vichAG/KaD6EL3mFwnHzfteunCBiO8X53iSVL1DN6w91ZB4XtebCo4b0hq5wn5DMZmTwzTKaA
Xq66qq3U0Do1cSJxxIPupGa/1YSYf4+McJ6HQdrpel3nnFO66NAgRAi8VE343gCNvBNHBx1X2psY
+auRxAMHaGVlgNuf6ZW2LE4DDpL+cZQmSgh7RrsZLZcQCt6XMRzi1cDjd5HRRcOD31GYDonOLuQP
LLHRWC0vxDfEvnaOSNLUUp7lj04/aH4ZsSPq2M9xgI5hNoOHf6XeXcfV0pWadW2ObmBbNZoITQfg
Dg7NF5KP6ItC/noQP3of6YUGFZzkMfRPokyF2aadII7UidM8kRrP2jsrSO3qyvlaq7wIvGXWZpuM
igV+xsuTI7rbkF1K+YIUXbd0bYoaD45r883lKYghUeINVibRQh43MveD1faPxqHMxJUNm34Z5r/w
9UkOgWH6z8JZyHD1/LHiaAnrSzahOWTZ6fpGIjxgBT0WiJKDAh9TWlzWZztsDmwOvwq4wtxfFhm2
C5LmfJ88GyqrYFzqZ1Wrw3ItUUR0XM3kh6NsQ/CEjiFvguIunnZKwsYNii4enhheggtTdtQfxgMN
dsJcFpsVou4M4RIm2XSMOYbGDjoJIMP5MWaCugNUaCwCQpyQXp9b6fhNrAY3dG1lP7LPns16b7cm
nw5wCeD8zfnAHF95t9gBBs3/q2qYYSSwutVyyyiotKCbXfCYHuLEgCB1UDaqXHHvXZlSJObpiLPt
u+GqtIlU8gPnFeutURQjLR211l79m8jveowKmbk4jwcsG4xYECABk64kIFVraLD3KplbqPMvyw9J
hXaN7QIGk9vZ6TMWV6nMiBXWuoR0QT5LxNBYf4uMJ0ahObFYO74jmNgIzJLQ9GpyS5XBWFBs8O+X
BFrFUS2mdLDR3im8CYK6Dcgd2xM3dtzYga0nBh034708dFe/IiPY/3a5620RcbciRfn+WmfA7o6G
+C8h81qfeURLP6oljpPcFNNsakLCpyumpE3strxp4XFdBb5SXgVbyKSBbAIn/rPWQRDsRDzfkqzv
YuoNDHt0gpzsQ26OmuSOj5CxrrA0YLVad2uTOmf3Fj6Tb1xN5P2X1F6Y4445Sw4P7ctm1zUVbW2L
/Mx6ECpoyD0ToYFnLPU4tC4DfKjkyK1rUX/oPmg02DjBVQ9bNXw9wxORCXkb4xD4pDvsU3W3cDpE
lRJbNRbJokJ58lTPLGTwrvkoIWHWEIy+ACZEyB1ltk7+fToW+IP528OATyKyjo4YSPqC1hWVxCfK
jdOTB1dztiSDL98pIKA0WK7v7joMjf2PFgOT0PDG4f95UdTsDO3KjJ39zWdg9LIHiiBJyA2Fxysa
2FqhDNd8GM7z3CVKHo7auXVDlVDPd4lBrgv+GqIHNiwMYybakcjpXDIMsaGzLywA5z/C7IEk3+I+
nJTUJQJQAtqUACl5f7eplOno3A9x19k//bSoorG1o5R9x0vS2izFVOUdfXXPuiDDWI88VVeO4oYy
h48JGWxazEACj9ana6bOk1rwqAUCMCd0c0YMrWw/pek7sg8IyiqTFj+LYxG/qdtAk9pFTJ45+M/w
6ReR/LIP7uo49PkYRgV/tthrypCbM9+ShikpbCul8btxXQnAW2O3908KDGhu4TkbzUIrfsgwZQnH
yN9+9Jaizh43igvlW4pWBHcbHO0vGsZx06SInZlnB7qjBvqIXKrWbY2O8FZd4bwt9zD6K1Wh8bp5
3lPZAf96JygqIKvBcjYIG9qwPINQ3M1t2ntrRMcGBQTZJaD0Z32pgeK1N25Zq6aV515ynCZ8ujbz
y9yKc1MczuA/nR80oKhfKUi/K/vNIfBgt00sPR6ne+ACi8NpVB+8JaTZpFkkWQ52aWeqM3hiZgLI
Mqk5FibGJY4BT1W09WpGDfhVwiDyFDAweymlLBcCTLr1seZMg129dl2XoGMGAx8r8He76791RnKi
ikRQWabTokjcplFUHeLpsRh6PKuYVzizR46Z1QzahYQll3cwciOJPs0HFe69JVFOm5ufR2NdTaRN
3DeeO4ZaQUYb23jFiqfSDYLXs7HdEqis6ekyjhNAHIUeMyXjvRtdEf9uB9ZmiI65HGxBx546p8XP
O4tTBKs7jeElZKO2qMA2lh110WpsxYj3rFCBY8CfUfV54KdWX+oOL4VjvFAHcKK1V41+78Ggsh2R
1JskfPuW547rUetcXl4/cCep66fs70Nd5wr5xAcyYNurjxvFTG0c33WKyfcR285Zc9Z4dlOA+blD
30ImvHCpMFbAh5iJhQ6XLr40QWPxuK0NsHEAiz4GlkNdR0fRvouLB8hKSMBjiyjB2JohMjZefil1
r7dGibyLGAMqXqs6nj6GA87i20GfM7mPhHtXDhFqr490Z/AWkZZ0uJmLuLvxiUpOEm+fQDv1o79C
HLhKpu+lD8u2kLEgTpj3NPvJTZTlzR9GcBUz582yu5VIRaAdHbVKQK24SnEuxPtVQDyC2xAnHr5r
gEtFeYwoGO1rkqWChhgYXXe0Sdi8ZlYmZCwzh+o6fXHy8NZhHmxXfhdSi2HsMA69MSw251pzQuOe
Y0FRzwU6XH/+nWoo0bfaIm1RJCoNgS631vj/YtQ1qT2f6NM6rrKQN8VHQ1yv5xXUr1O/ZPeD+fVc
8QTBlCJ9NtiKOTdMG8xbJC0i+WllGWk615mwNuc6Fng7LoM8BXfzGw3gEygbPWhAXT0mVCLzIbdZ
unI58jluuAd7kd0CYg53ejwV70MBjQ1RKWgS/OxN8jfBhgeDFEOKVYeUUhp4Bl0UdFLJO+ztLrm4
WDdtIbZoSiujgnX7OLp5fgX4PT8J2sixQ2GZGAJ2Ch15fJo3n0cc2M/cgP8x7A6gGBUqhPpeEw7G
UWaQZ2YL/jE/z8C5QJSZQ/IUVNGoe3i91oqU3DUid1OSwmTIpQcN8b/JR/QEt2zcCC21joj2mh8p
mn4ode/82AVNLOp2LSkIzqAeIH+7Yku4hXthRuQEPWjcs2zY2/uHNVK4/H7g87YuuS9/fUpaYbwi
DrDu1+MWOi2Nk4sicT0LSxaXtxUT4bd2eW5cQDwt0cZit8KmtqNtlH0li8Lm1EzkFBXD7LpbcYea
OnX9ZzPG5Cah1wYT5TRLBC5h1BhpOv2aXrASBxI6sEmd9Cnuqt2CA7o9WtxWCz1LyE+hkExVZQlY
F4og8hD8jgv2mj0Ngd8EmGbUfh3ijAdd0hlYVShNzZUgKDesJagppqzJkAgCZx+Mhbw3cYV9CAPh
0tLQONY4AYT6dCEFifOXJoufajRLlOw1f4jCxH0+6EsEKkcgOD1u7oKhxyJmgiePwfeK/nhfDnAt
LRzN8vndViBqlzJ3USLLmeMdSEYzbr6RHJzRqAmTuNdlbZJmv6zrUngcfKRQreyL0fTBIrTrYDxJ
2YLbumMR6FiV7WpytKzKv/mChBvkrhAASS8OVMllffivmsNC+T7uGWPw6aXiVQJ3mukyB5aXgXQ0
AU40EmCaI3btVdiGNT2lYE4Go9iho0kO45OYzscOP1PePBQ2DXWFSRSyZPfquXhkmaSGbMDW7oky
J2P3mtWlRzRsERaDN3j+HFg6bwP5emwassccAPmT8S3y5uuGubbkDfYQwFxbbFDXUR6BZTRUO86s
S7offnmbOi8DlQflIiA9ZaEXqfykVYT8/CjwoWoDB+hogoLT5TqzdzJAzQGupMsEJ+wnFEVnXkjD
IpmGwt6FI8ftdJeKcJJt6AIdQoCenkggJnqm90C4I/TlOVZhPMLIS9hb2p/qdevqmjW8jg87Y0hH
vnd0T69vk7oXm1emW/XCNtUESWhk/qFEm9tj/61B+X7OoMBTOFCzSWEBTBysIBKGYGBJUGd1pA6b
UDTXaC+AiHIDPGURito7Hv3vaqqLc0Cm12sI9Y2DgDLti5ltQ0XsSAfyCPomxIFGew0yVDeh28lo
58fEcyXve5+yeKMd3Z9m32ltLtMJqxsCuSVZA4V2Yfz5y7a9NixMRqsOHW9EPmAyVouS8mkp2E/Q
XNg83/FuJV6XzGjF2QUY6KPdsWfL7WbgaYGQyM6g3GEvnZnyHJw/Mc54su9Cd7c/xc28fX+m0Y2n
D/rhOdFJ+tRq7410Ir8FOk0fmjMD/3o/oY3AHHz+8wtJm5FDL3qTz4m5LusSaBAkBGoOlYvSZoRe
anNNDKV//HE/R022r2whMfHj30DT9k/Vu9mBEmcEVBUx4nP6/3E8I5fjtQSdBuPDbFEbiQAaiDU9
l60XcNqJUKbayg56XIVjhmOobyoYSpbMsb0jrDWRUr7HpLao29tte/bHkcxgI2BJDVlZ4KILqhZi
iDqMnLpffVXOryKl6H8dHFxJFSixO4WvX7UsfRPFzT9d4F9uxd49eRBLIsym0vQlwDpoDo0RP4lK
ebYzpOr45W9qmjhHbrjCFSzew1RHBPhxmlYzB7YoxA8jfGNSDitWTz3MK06v4e8nG3343In7ijTo
6MuYFiqSaYvmzlB9mAnHThPKQVWooFD7FROuZHYNKLDQX/3W/5fHQbL3GDbnn+An0QQN5mTwJfDk
gQwdgxo6kxi9rLe6fwkuebooZwYjud4nOGW6ej1PPXWvK9U27G/rym0Pa7hwqPdHPjMkzDKhcRPy
kkSbWJfJJHvHlsJyMSFxf/gpwV2tyE1nX2ZFcrPVMCkHzsXTdF4aN76A+bQECqJxT6SJ+Z8kG1Uy
mDC89im2SlrjLTg3Q01EGummu9GUYiAu4BxBG0IpBOpc8sYI7dIZzRj0/crZSl8M7Zh6/ganNhDV
3U/9a1KhVH9c0wWhhNKxeiOZ3n2718Tfd9WUk2fzH/+mSQBZmGHb1Wa3IgK80rV2r7wOzzfYGHHs
NFbNtakfP1xjl8B4vg4pgk30RqBTDSi0ewG6CHZstAsGM90TozbY6pibvjE7FtLRPbut5AmrFjmc
nlfmrbT1sM7hXcGfT02lxQYQtsdoejPimWEZBPkDa+1YZrO7ZFuv8qzE2xmbsUP/iP9lg1odaAL3
q06kh66H7dD8IJhtmnCR79gH9LfLJZB6NaOjNUlGAtauMa/98sNdM3vBr0xpVon/yq/rvCv2qCwD
BmvOEuZEH17csqRsVJj6U3x0gQmR+xrbk4rlvAh1kJOkr+NYfxyrn8eFNydjWJUW+4IlZzKLfBKI
CIeWyAQikiSp6PfPqXF2WR3FI39d+Wl+mKhk3HHTzsnzgODP3BQRTyLhjREeZFhQO70k1QD0GPK3
QTLtudv8cd4bJxIvHNOF0dqReDMQjfx2UaaKlG5uKtC5HKY8QeXDdmxAjyyVM6kXv/x9VccZYzVB
ZtzMHRS2mcrlC+z5D9bltf5OrPj5UMgUWXNgiRWauOb1TtZqQ24cobwpkWyW7Bi0tdb9uafBWwoZ
GD6Khleu97+244v+mbzXpMNe9QdwBjbZLavVbFHYcKHJA3HdBP1COTmi1iAgtaemnckSR2OjFTz1
adKh4wEro/fs+qCITBDDT5BXEnZT0fhWEvvxfj/PFMH6P4GbzsJ1WMWF8IjDCmDaCpAgy9fOF8G6
xJTIQuP8HZLsfrqzR8Oco7r3AVmOGtC6EWtmwkWJM1OPd1JQlQC9shEnxvke4RDvJE+lVqavftn/
Z1YlmkmLmvoEtb5+4Y2OP/pm36F3rqIen93Gs26DrQU7pcCJ1acNGRkov3+aVuzguaQ4sSj/OWcC
yM2BYNt/L9wVrZ9ZrjP15BCUhDkcFAxx/UxJWxsmevg1Axhkfg/OhXR82h7zDlPeR96kVAK4/AL4
WZV6CKuSttsV87Aqoo1dDw84KaafhWlTntPUe1+OYpoZMxv3mjU+ebgI3Lr51/dyh0TrbV8lT2Zy
ySTL9pa+7wzhL9nGxeM98lzxLQ+ITuuTtoLaYhIsotGDHd780x/qcCbX55nWmHqMh+JBcEuvaIIm
+T0YZxWi3HyrR7jfG0rkBGelBxBz/NODusZESKZgNZbNNkMbFvfj7xNCrwQQHEPxjhHtEvxJ/yn4
tEFmZHxcuaXNp/B9Zii7Ar2GnwRqdzoQnP85mAMXtul7hYsfqv0yzR+8wQ2VfdzU2QfuiNNGQcvd
36024gSsvNcX/217k/80GcIw28vB+oIaidPYa4ofQWPE/xIEYD2OIXR2c2jpzVU+W540wGJ4rcVb
wCAIUA5Im+xOMG38cq2lKh37rsnvterxZwY69BhqG+Z7oToAvyuGC9G5woe2RrPvm463RE/ZL+CZ
PHv9WJqmGHwNHRNGbsY8C6O6rL1q80GWKeXwQc252F2K2SrHAiAE7CklQxgOlkmYpDb/ALMnrEri
Y07cTWgYzEsLFsuUkNjDDu7fr6MXxampI1VjekuZj4ewfrtXvahXUjc/+6mwXhwM5DnGAeMKVAnX
pnPLCbCXe5l5oiKSAPi5FuTtoRka0N4bfJFo/1LlRlwC0tz38d8kMovqFWeH4DU/0dfaFXPXQ9Ev
PG7RVDDDxjbZ1tdgpxiHrpos+8Y1qP1iloCiECYpXg8CyjTjrsBokv0sm07KMJCjuoBMgE+93U/e
EYYHfBsiI/6o6Ni6Xy372SN6Z0NqbluF4e8xaxHY28YrkdKBXOeLgv0ws1H6uIQ5rBl6D3mhwDnE
e8mrBCrKNSN+eWDK9WMJ6dlDiPJPkpAZL69yk0RsY+5H0uISM7BUyyUO9NA2CanP0h5xdD96lAHw
1eI4xm2wp050hVdi4UbmpG+0jZAqvHA/YpFKLsaOb4pKl+PaPaX97dLQwIdsVtALSWckmj2EFM8R
T9rtyKKz45jgS8nTo+aL6IEisF4qkhqR+sleb/Htn4gV56zOmkqcFO3Qa+8cjzt3uhiFjPd3qJey
jsC8UieZS3t8Z3LgfoaTEtDKG/TcUycHD9ZFPMcwnKW5dnU3hocCptj7UrPjxe1T9V088dcmkqRe
/Trdjv+6QCHX5t6jNX+FYBBT2J6dPpDvLqtSPAGPz0AWWpcn+WqhrptlKNXjZ1LuxThJruU90D1I
No3N5QKFrazKJjNtVkXlvciGMspbwN1lccAFbaKOOd+i9MYYC0j/yaaeSyNn5MeF4L/hmrCY/HoP
5nAiQXn1XEjYsP5eluPZIg5U13pS/NEoH8T9iHA9bpvNK0/fdZz259Snoq9cGyaJVHjP8LGBD+fv
y9T0peIbDp6mBjtn0Hhcsrq1obINApJvTEOlFCjo8gNOUDkz12hp/uVrnIGksCbUn3BpNtrrLMlv
863qhIB1xlfHTEMYtw/3zi1FlZ0O4W4HIInJXgFrwa5p4G6GxW1fdTSbvUjMy0JmAe9zZ23gCnQP
ycWy9NvO4dwauZYtdNLzGhQdhq9sCL8LxKgQLjDtDu/FFHhqkCmkg6C0NEAmqQ8MCzisUDaJ/rKa
vEev0jByIxDSyU/507QX/DFevd2cdTa/L7wqgoYJlPBOeqFbZy1PY1L4ud9Nw5q1RpYnDl+iF0Qj
dOrhkmSWxDHqNRKqynWfvS5d7stB1I07Fz7WttwF0Qh7/FggV0CP5CeAA2O+JO/iscLWbe1un2Pw
lkwbf5byzCmEqyMxeFYg82ojqKuaRmNqf4FLNC5eNAWLBv60dVQlDIBaLHuREmXVRRfmCKaPmxiF
26OruIEDCUur8In+IlcJljRhXGMaL61iS7v3xqRrMGkssCxq/r9zy+yZDOaCLdBl21gB2vFR+xjb
4BWki9XlEkdUvNkp4Dkd3kTb/y0nr6qip+VvPQIQQVYUjaQUMBfwRwC1YKB/wXo2XETF5P3ywZfr
ScaFkvix2Upuie9J0Jc/1SO2nlKVfUCEs38kVLN/eYULmlfQ13Hs1YvWq0C2LSKuNK8HRq7RtGC1
F5IFOdBcRMtEHbAxOK2yc87YtpDyIKJFgItWaXoq+UdTN+IHgTqJrkhEhaIxOSIH8XmFm+YqeBuJ
TSXne29+xB4rE5uOAbBKuI2lC7XpON/BloJKLkxqJ4owb5LZ0sqfEgtBIvl6oFnciGFw7CIZa13Q
61EYngQpuWpyEFMvVHWEXUfYmH8pTWh6omxiEDKyBhL4rpNndAZX57ngRZtSQCSwaGfv/obJgx+J
NdT2DZAfOtbFR6WmZtC/B6mtjg+H1kPb5JAjLCjlBAJwDZE38E0rkK8q3fpNqFKba0L+cN6+fPrU
gtrBS4HPyWm2XCr/dLfDYNx3d37HLZjLS8QOt9BnYZ0RMq/L0ae8/mJz8rTRcghJPflcOlivdEbE
kZ8Q/VAT29V4aQ1joE3gNprvDCcxLI4GX7VKkS/FLdDgTwiA8zXMc7cJGlxJpOwcDkzlAnSFxHIk
KTapdQYhRe8bvmA2fz+apegNbM1Yrh4A2a+40uhBjjNs0bRPqJc27WAuDLfM2PpJdqEEgdMZYE10
JfVNK0ImjOgbURbVYygPBRkovI/p44paqND4Y0mv64fgq2YjJlGXqzui5G4QxUvBK8bA1OasCUUz
1jshgb13s3PyVvlk3pTb2iRR6B0nwEDBt0rh4xI43ZH8az94sFTAb2yBFfyPgWDGRd/NF6UrD9jT
cdyFymnVg4KM9F5sv+7ayiH+WKLbZ/FwVSh06os7aBo0+YTL2MaL4UngRU3xfqh5PsKLgsu5isQF
b2CE1CD24Fxkot6r7Eu3f5/CDnLyudH9bGvMsjbFAkpY77Jr3KmYsvtDSZrxoeaJA67WU7kBcAw1
INefY37LDq1Gq99WU4gV75WEqwgj25UKKZx4kYrPTapG+C1XlPjlFY2sQ4msMINZyOwwJIfz7JzQ
ydf6WrQzrIMhrfa0aK3ImCxJaglMxu3Ai0SFVlAFrWbr6c4GdkskFZW12wzeRGV2xUPO4qvhMQFM
hg6SgqyUiVkaJf97zVdS/CZn/nFUvSUgMycOUZS/vPxLrz7faFppQ1Dqie9IppUBJRjwR7e7c+5Q
OEyvlu8Lz8vXr5SdvKpFeji9tH1SRASITTjt/y/J85gHGBunPOtxkdOZ9CdGw4EQNJwg7n/Dx2dB
LSjrMkvpXbY2t7ci5oVXnypWx0rtFVt8GYpb0YDDY1UHND91C4pWAH/qN6/tabI+XyDKxjoyJ6fH
WeigwLlVxSYqU0sbO/IvGGH2PfN7t2M1ch7txo18P8GwHgsgj6LuyjQo1Kbg5EK+FO2Dwl/FE/jD
ulEzRMJM8qjrY4jWf8JhafEJwc4AcSdv9hVzIdms2RAR8LIMdbYh8SVtm8guH1e6V+cBB4K/Q53i
ttUBJ7YFAZLpIHd5LrqCOgjjKAWIgoQXj22puo/OOcnUZ7iK9sJPOrb8KQITzjB+iY6VHoPVoM62
7u+Knk7scZFAezN3Z+AFHEMjFmQStZXrNJrlXwkmP1E/bel8c2Ibr0EICMCQ9rv84zTAbkLkgUYp
S2DvwuFiUFM6/QHH+NhJN6XSvmMDR/lhNLZy2tRediw1Ao/PloQtXbXrs8qQ147Bs1YD55EDwm5a
CfrfsLmYm+ufll/LnDqqdahN7A8oPbXTOpOnpDJG+qf5cZ9WKQHkqVbl13UP7xQohf42gL8Qp9SM
uRuMby7qn/Hq/+0IVZ5+IH2fQJQxo8bkXaFZuybJMU9ew9BPbRaWbzAGWYTX2iGZo3cASUqQUSny
J5TRWBo2cux4/Qyv9ce4L81qlJ9btYY+0+nBHkJVOkAzrZTg0GD7Ar39t9Je4S+b5rAwP+3SflfX
ZoYwUG33kT6Sk2iMLq9sePgF9W3lY9oVdlxEP6MHQf6w5aT2DZPNvykU4DN3sIrZNdNxlbiW1+6x
NrCro8S8U73zDuVsjqz36F68p/OyQecLUm5yLmnIdLn1gKlSTDiVQuDeOpC2tvaT6L06AKN8TK0l
M6R40mOg6hY6dwIGnuNhFl3ICE8epSmkX4Nd47n7rErs3MONzQuWqwhpdf1745Bi/cf/nRnnEy6o
XdUIrN65h1vECm4312+IN0bx7D0Ky0v7P/jOwNjUnnrxC6WY2TGEw8b2rX8Wobf+si1VLVTDlgO4
n3T6UK45OKWbunzPN2LR63AOxaxAVTQezfaa3huo9WjBKutoSVK250V83VbKUikW09bhV1rZtQOD
NpUPKjlI446qD9vYtLbn3RiMoIFUbB2mtgv56bjHAFUV+mfQaXf22jBHjSodItAKMb8LILEihGAQ
ltP2nkXezoBFXsUfnObvpRcPf4tnAH5ZV24g4x18cvm1y/b62DkltdAy3MLPqdRNmb6AqSUWN/Iw
C4nPvJ0RSHtwbwkcLaCb4I8IRqM9bNzDMjkTTUKw988Mr4S6DYY25YgflvDx3kWxWwYf98PiiHBQ
dt3N0no8DARr23WZ/g7Lk/Cw+juKYeIMxLpBN2oQNp+0Nc67oiLqY0IYKPzn8gPm1V5TICdJYyP8
u3swUYs6YSbf56BSdD8Bh6zqxpLi1P74LHDk+mYexrU6Lws1m58g12bbPwTa+axnbCWCDwNKn4av
kKi9GkvV6IAUgYb9oTonZZNq1qYB7OMSYS0G4YRL3AChs8CLKwl16oAd3aT/vV9z7V8S39IX4sjM
SOXi9KxYVoQnFbmlIK9oWHW+4QII+A7lO9U34yV1I4jD2do1bGgPh5ZdETnckZNuDvYJTZew5U42
SLP2dhLNOK1NtqyE0BVRZRSiCVa999HWNxEE6dPF/fMN1vccPs+lhNsCp6qlEMgftBsBessdcLM2
mxZzcQ1cS1Oz2Mc5QlRbh0eElKUQeD7p987k0znqj1uEUyi8E7api+Nx+I03Y/mW+nu5jP/MrKXZ
6dY9RNH4+0Sc9I0P3AiWPsgC7QaHCZFqiCRzpXgej4rhPUAK+icBbpReO1hjYDZ2blfnjg7aY2bL
0CE8KFiFyVNQiwRfYDMjs1blNxpDBBxu6YB/GY78ftd0UwuXJk2ffQOlrhghZ4c5p3c82rDyLT/n
+Kg9L8SSwdIHQbsU5f1zyWIu/UTQ6N3DFgl1+5ibyZgf+Wa79kSWzw3pw3NlGrNaAaDb9ocj6Q47
Wh5igIigKCeCdp//KmuIJMc59QQOxU2ncClHFble+z308W37tHl5wnbjhs946cRj7bPgmwF3cBdP
KbaKopIDeys8ew3yTlykIHcdTREkfj4D7pPluuzTZUFg11F+gWgl/rJbS2jy0w8VQYY64O70Iw4d
6OV7ScVrkYw6BZfh9H4RDpRtR8JOS0QhXWd18DdLGpyrDLTRy6Ful+kTXhIgHdbJ+wKOds2eUf1m
KyEf4zHI2bnOzEEg/FlcmvUDMAdg8u81H84gp9Q+LiiOqtcgkHnL9QE8Fw0/YAMPn2IkOSBuZdFz
oV1+pAD6T49/cS7OC3x6sy1mfTOLIuc8VvPxuyM2ZeJ2vnuM+4xfBbj6ODuTsjPT0OyqRFGJo+3S
4X2gx1ahaQ1jXtAJUct2jWOdgyPug66/f5Mbw0i1hMZAfxVnnGX2WADo3QP8bYhhPx0FepmQjg47
pmPfgPOU0nZSSrlu0GBtyfT2gaYiExze0u4TirVC1WpBTdsF815phrqOpDfraUtBnDWRPYLpuqow
nd8/P4SOe7Fd07pUUdFIG8n9H4IcdiH5kJIcYghXCbTKbRj2VRAQ49n5PXvco0QU2RlLjYn57kwM
mSL3i1Hsx2lbwqy2t1X/8u5c/2uumkT98KqZfDiFPSMk7/y3c8FFhXEmkc/C66k5HJheqlyrNXH9
O8hSrDh6RetRagPCyOq+8z2GxEjlwe13NbRcISb0xEDKsWFTKRhSHH2AqT1QHKnB14uCMsngX86p
aptcpSsBcIclUk+acpEW49SG4wbXKtlvsb4grRxBAtovUiRX0f5EqeZHppqspqVEsgxG5JqXHBQp
PKW/cuj6T9LiFEAXETcny0V/gIQ0W/2GN3R2XkSyb6+gRduiVOm0nxE/srOnuZiwISBslo1aVMYe
DfEnNMXhcbEI/wAlJJ6LTZkwtq+N2yFf2+Xr5bVEQQQ2ckGXyeF10AjeVs6lI+wQOfDeWSjr1LjD
3IqUUd5qDBZPBzP1fq6u6ngGGOMu2zzOYoS+VNYCfLSJLK2H+rJdM3zaM7k8DPdGr4c+smlmLjtI
6RC9EBv4LiGZiGzKvEwFWvp+ctVDDHjihPqHbvGGxkhwiwnQo0hiG97TSTm70mWK8ST05xsRDDCE
EL09jzPHu0ElegVco+OaWcFT2sR4MGFMtjZB2N6ynaIHP4f0UVIPL1vlwwHa2wD8OOs3ZNSJqfKH
wQFGEgHw+9//WmJiD6ysrHImOh4WvUDr8JMeKFKEuKnRHXrJEH7Pf9NjdYnT574xmKgEGgbWlgFn
CRVftO7JtdDvDzXjGq943Ti4GTE+jhGa82FVpBx28+FjwMWJD7B+mmh48NmiY8lGgudCRDObAFno
i87M5rEu/hIE9E7LkQPE5vixIxf7J+KXY/9sadNmzDJUGJ8KkCrs8BfBvnHynegOquddJmJFuIwy
F4YpYr1W48KDGL2pXb6xVyAbeQ4Fja+X4SxZi2eBmsa6qugbTcVBujRpHDXvJgLa7jekNzXBnDfl
Xwe9YCq1dT6PvcQfzGNyK6+HKfSXRZPoQ9uvSxftl7jHr3M7QLk43FntFYkiyWPug1Elc54Nt+6z
Y27JVkVS7avvJ8Cuk4imxQeBeYDPs8DARNmVKOfj8xMblqnYXhxZ+5mTuv+MA2JyZH2g4Q2whdbo
sVOZ7K+EnylygjFPUfDZynDr+xW1msUhOMzmazqBJxG7qmIuSZHMKXht9uMfzeS1WCrFd2lAF69z
TjpcfUwlOHKEknHgQArdQfpvw0rlWasb5kLSIioQOX0lLOh5VHOrPCyexCLwFSqmxTaoeNEPFlOb
hgpZ5RVx/xd3NBUgr+u3Vwg2OHk4XGrk4L9HSdmFNA5KRIlbdijTqx/b/jmLPye60p3tzZc2ckR6
HL38gVL4n2dQt/TWjrtWiGGPbD3YucHtZzedKlcHyr0i4bfKwZkRCvDWAItoZFtv8IMDOKd35arn
AKC1XPeLr4B9NCUoavMd/asIwvnI68mILUtCjV3LGfgmUjd8HjiK5XiQPrmogjnOUw1Oey7uj1GV
/daL4aQpVCK2Il6Cx8K79M6P7y4mbmDFXUBVeB4PRHnVIZZM6YXikc501qIPyn0M7ElbdlcPXG3A
x2Y3gCOWM5wUxAO+hiN17CW/cNF8KfVUEjn4s/W7Cd20Yu517dNRaU29zhEORdGK7F+Ab1N9JVOS
8u7ljjklAYlGE10nGvp6aJ/gS4LNydwqqEp67Os2LCgidSmn3t/l2xJeT+qUv4Dg+RlYiIN/sipf
xIJV+jxuaWzli5BkKUE8LPkVqEiStvi7ejz9ZLkSFJahMCX3ZTusnpd0tQXRF+Iw0r2+2NV53zL+
qWwCsFX/EhjeuLQrrn3KAz8+LWedoQBXVkRaQgkD5vQH6FQimiswXv0lDaF11yZ5YMfIUQETpcYx
irRAj3nP1iR/WCrHYDtsW4pP3Zken2mujFuyG5Him7+Q3KCSeWeKwD7+a2YTMyh1DDtC9DZ8/Unf
J/aaBUmtx35KzhvxvI9qyTQsaUgtFIl3wKA+97tIwOC+cyLSZaVC1CRCxjnBk15fSnboGez0wgrg
0NQrm41SoQLEw7wZyWO8q89dgxzmMe3DI0zZTBE6fbrHqXD1xt3KE4SbsyvN5X/HcMKkFOgCNycp
oZYZ5oU6h239/9Zg7j/rh2TwaFErTIv2OxMlPajrO9KjGyYCHvwQvY70mZiGYp3mB1aAC0JS8wkm
lwdI9ph9yyL0FGDH4zOBM9Y++slcNs9XclYdE1D/ydaiemBxZrCcZpZO6jMNeO/tVNXVcHHsPleU
MMzuupMDxiVfEHP7+o0nO9TqdyrRjJyla7OdwUOZdmoTcKmJOo3u4l2+6QBCwLIIc/kyq+SSMgpw
b5oUziszeH5Qvcb7AQuQNcJu6YJITCuvIlt1eVFQ9bAR7Y1S378cHkWKmzadTqhy2tE615XAbt+e
4xd2B9Sw+85eWZByH/ytq9FCXxTtYzja8SrFBjDDjaIJww5voLHyx5/5cVbjJCSMV7HkJE3AifQW
5GRMKtjB/8tiz7PV3l0ISXV6W4/WK/UsVxFjgScO2eS+pymUVnsYseutVtNAusMCMFT4ZixIANBZ
WgIXc4jqRT+yuCvZcjzbMB0FbrwHa+bFA1Ob5Gywefs96iEEAoc7MlK5CvPgSrzsyOiHSowbGKVc
l0uOVU98xCAPk3FtDsh7BZ9j+vnukWkeLnT3FgfHxFOM0sTFAU55Js7kkAY2jLn+NUWizpx8e8fG
SUai9W6TbTXw3jRPUDk8gFbVgxZ+oJJl8cudw8UEvCu+WO1ytanqPnSWHJjWLKkcr23ggqqikgep
IBxELvlxSzCgBzTCB1ti7WIWY7IZY1O+w+NE9J1IhxvMLBmDoOGbf0lbNpCi0X36+TQ2pLM1qupa
NNx0dxOgn+fvKqWadPo7UCvFVs+R31mVQtr4j4ZHXLQEoRFKAdEDqTeS4M5/BHaCq7SOqk0lCtAF
L4UT/E+XlinHALTJrn97QXnNn6vZptIDBPlJdXlNTiqgZIGN+7FVeCq61VrDJMfHK217kLA1by78
z2Cvm8oTXZPCIU+u8iQnm8KxEfRd+/UXs7F5zZPYfgbLP7zFatooCUBp9jYIazGJJ0l3XmdZGDGF
lmEoAhVM38+bkVPA0dOja/tZjqwZqJKYfTmupPrpO6sxdz5+tT3/zPZgePFd4ulu0MtAKvxwON4Z
syh+J1h/A06vIQjIYv94pq6L6Eis32P0yDbT+ht74f8hmgYooPsoFlpzfZO4PrBTj/lWedI5mf5R
fE+IoTidMEKJJcRXkwDnFmb1/ROif2I1d126LGvOn3en4cqgQ6MVw149M/7qjnz2kHWsRt2Rk3ao
85dAGhQ0N5UwVyC2gnBMdjti4IdmJ6M6v82wpwPAfe0If3wFq0ADYIMj32sqL6oIwa8Ibk9+VnF9
NZqWPCmvq9DbdJmWNw8SAYxH4SsjzV7nuYUxMezOPiFe9BIIGl5fu+dBhaU0J9ahd1syyr87cgQo
tY3zz3vH1k4juJysG7Dn6isrci5FPDHXtAeKRtQW+no1bau3K1gzYmP83nhzlPwG6B6AX9Nx0Y5n
NOgCxAHKzT25ostjikPb9a2TxA2TwHlp6SK3pPtjq8/GTyNe5s5gIBCnRS1ESgri3vs2XnN2or5j
shnKj03jmLXPGTuNkP6lXMSfH31czFWNW8CJS5B1lr9AA1LESaRyqpTjgiktzhDDLw5+goSV/2HZ
1iDtscfewb4jPXZIZ8m2RCeOm8oxQqJcnULt1YWq4U5MOhuIgjV5zgOThIj7x7TW8qaBd+fsknQh
WkErqOuSskzzB+ZuzgguL5wVAQ4iJn4PCTAnXORzHCfWCaZyu5WmqxsOux/mMeiA5lDe81GK77y7
QcxUAqsqMd82Li1ADnUXznz23QWPUhUt7TPffbCJVZEPb4IgsIlgtQd2DLV8OWjg5MZNh9qh5PM4
HI+PHCAyBAizfsz9yJ69O5wwJWfBLNNxGdQP8BjYNnKTasiHiPTU/VcIuezT91i+aM37G63pflH2
Ztc6+yx+0XHLwz19GSxnWsNwX/oienIhXiJJqbZz4T6hrVfndZqATG/OzbT5wogVgTm+GzFdwkVB
X8ryShb30FpNSXT8HS7Jtv63LxbOFamFhlpg8QJNqWqY1NZSzwhbdkww/D6S5wKAGNMCYlyMaL+r
nwy2xqAkM7j57ls1un8S/09XHGUhm4rcUaQW/2nyoYe7Y2dbiDbPFgcLGrnC6iIj2qMTpWALerBH
a79VlXyCh6+K74i+lMMMDgzZZtm0Z96aaJvSz7N7AUWX6Ybwo866c8z2vQ2qImsXIbZDI9onww1R
q/pTFnD2ai04DypzIOptAyYbQydgX6nCQgBmdbCb95A1eJvAkG9K3SEekXZFBrnD40E8NQisdOly
ndRcWhiML3l088AQO6SEQxopmdYxp6db5yDM7Sse+ZJwKKk0D+fcZkG1P1IaxUJ0k43TYIGzXXm2
+1fpMU04UE+q/TNfw0jIYqEeq8ktAQLW78sk4LoZ49FcnmflxQopC/MmvkzD+9luO1+21ZpENaUX
8G61euDC9wAsM75/knwq1A/nUndka1RiWzvVgI8usFe+8XyPHo63MWl8oubJmaFysn1WkkbWmofn
10qAdNAZyNCVeJoZhPZcjbjMhuAx2PAqs8GbOCA6GXTb/wcnaAcP/aHqdVZCzG4iP8ze4cFGPyKN
PB1Dm4oxBkbVwlO8Db772aCeyyuBxhcByRDU2LAF2hmfIf1KmZt6e7COKHXJNeW7aN4CKdptY7aH
z6+Z2UGF3yxxKNedCSdPQDB4z7gwAmRghPlHNpxlAzWs4FnviYzvVtdj7mlHosqvM9PcK+jDL5oO
HUEPUW9MARhTOZaz/b5hz5e12u/Mlvghoc/qr1NoVgbYDpQKYyqatPyhdimaiWUzxKZUaDTAa3sa
FSM2ZRaa1laFln+bjhq0scW7Mlirkp8rXjkXex0Sp7oROrTUPIQFTqz2zTbEA8SgOVd+gCYtqEFQ
18gHgv7H9w6lPVnc6vljAk+hrzRJ/uXTugrwN38sxgs7UdITUOpWywBLhr82Ln2UBvIR58v++IJj
Zw/EUDb/T2u8jGBFguJfyJcRCwipao7MpRhTvhUSgN+CG6JHEjUd5MzXtgP9VrFiKl66mb44YuEj
aCQdWEYkKCEJqp7Uu0QFINyU+zAvoc8XAV6luDjLSQV9zFql0D2ZohhZTfEX1teU/tT/LARzaMkw
w3tIR7fLu9VN/7j/0+BwmygnNU1OF4jXgf9F2TCRZ7VHPJcppmzRy34FXi14EZNwcaLYCo7ad2JH
W/p8/lNwuk+nhiZ0tWIHmtGedCzkkNiQdUaXp6OvmmEHXUPBaGvVNAEmnttYVyrAjavJ6dzV5MEZ
+Ks78wGm5UcRURONdvD0s/dopYNZS1EvZ1JGdsFmhVGK0hWklnc3U8qXfVjbJXwun2+Cy5kCQKlK
ONR+p54/FvMKGbygLvO05qCnwLMHth47G67Ez+RdSsSkyKgowUfyAa//FiCAOSGJA28QgedYDqbC
6wWS+dXm7DbNjjbPBKwPC6Mt7N++Jltn4JE7MslVyDwA+kUEiLLw30BSMtDujTWSWQQegy7GcRvq
62r7kmyCmOtxo4RdVwB/zaS1cHKlyuXiEEcVoi46aTarypZRkikWKNMVQcvSp+LpA6TMi2Qjg/ew
CVGIs1svGKODEPohxIsHKcJeTfjCnR882Ho27xL/g6CVJsT+BBlPtj/z5n1btoYeA9gpu77Isr3K
4tjWBaJ/Av9JAgF71nUGDIrjQLpHFqEWgaQdO5O3G9BQk7mpUqkROk1HQ8r7Ppkag7WDku1Pl16y
9I7B0RauV4tADhMrso0pcXSThHiHDZtcGj2QhkisQtIAD/J2SaYtyPk1qRzZkhQPP7fAp4kO8Mzd
QPSS4Ys6iU5PFksEj95kXQM+EdJoS7O95vinOeFU36fIf9Vh39SYL2sCSQoxy8JdRFYX1tpyHrS9
Y1EFxgdlo/5Mltge4YhygHeQAMoiT7tlbx4LmK1xjkXs0eVh2GTNWK0v9O9r26C/uKevy63WJ1vB
YTbRtkqkVNi3g0W9XrZ4HZbhFht4O2f8Pv6raRSWkCDT4hTi3SUZdc7ZfM2AkMO50EK1B9UvQN2G
37Ui84CnOy3t+21O+eYPuzuxjyTaxF+YGK9ZNou+MSypGPB24yxwJ0phzOchD1iRc/mxEx8Mg05W
S5IbB3SfbbV3adPbYgnc8pfXElJkSUW060/86JRtM8z/083SlMV4xj9GMMeNrkgq+6DMr0MbYCJ/
1Ydd/ESADJDpE5TafKgqBysR7wrb1nnivvJ6cCdsBEUXOhLG0wbKSdrzTWQJGGUPqYs8Y/5Mvozw
0BApHeYUy1BzDhgCyJFjPLNQL4Rlzg4wYX84+ieot/oH7HGZLUyC8dDj9APrsvDfhaEM3W1nBq4s
swa0cLbn1x8aedtw24oowPFS02fH5T0AalzQ+QyJJQZ+mQXe795HVnrodOyoL21BMJqWSoHYdEU1
PUSu+9CfQ10GOAi5DbfJdfibJNj9aDrDuN7PjzaVLUAFQzlseWxXnPXWhPT6v/wP5QA1zaGB2y1D
lHlo+ty6WwEFNpycPrlQlaKo67eCi8zDA53nDafgLFwrJNopIKDf72th6cLpGeXrfMoABblUEkAj
jtsbwVRiC1wFoYbaj/7bIahiXMXlkXoo/VtybONxGjlxA0UStaiI17OXoArFEeIn7yL7pqP/0n98
U1jmiX+l1uCkcY4js47PAmlJuhc8GzZH7EOLyp2PG7yP7BkZST7TOHKGbcuSeHAG03y7JsR5NPEr
Q8CB0w/G/dfwdAhlCDUSJvV4oxMe7yRI2V9TaW2KiAxP2H/pbgpRAqk+lEIolAFpXWz9tBJ6iv2E
NeUNDftiIiWQ8CyMtjnc94rn/xoyICumQ1vQNLJPZiiND5BmWFnzfV7TkQaN8b+EXT5R/CEP09/j
r1O1wlSRFAMfBxUSN2eDIpZdWc0li955FWr1KjOnAXvlHTqqfLxLpDdTZ+5cyv0WJBPECYZ3mq0S
PwrWpM332ak9fDuQNbABjcD35pOpMTx9ohct/b9vVdfCblCxJoNLHg9IFyTcpsjsNQneatLxaKhQ
WmP7t0cN/3awGBCfXW09+Irpexstcbf4L/AjhIP2/Rrd1n86co4ephafhSwf6ypCXecBRveKDdrj
jSInTMWMMiXn/3z4Lhibu9mSih5r8KyCoXYHGTa2sQy6rkpLEJMHn94/1Bt/rncuDxaq4dgr8Syk
LWKMBEqIq5Uz1G4MDSRfrDgEar07K/ylSKP2NMDe4QKrNutrsugckOV5znkgSTtYtyeTPJp2zsRP
5crg4Vii1hD4vOmxyHH+tTA6U8dWa49kW6Gid8JTST33k5TW8A4PMxSm6hbwTphlLrRoDtl+Bgst
9DEKixcvauDHW35UifSi01zquJmJ9uHxJlitqP+ZaRXoauSf1h+rQJHTYQ8pKi8fDQ+i9oiR9Pms
chR/aBcPwhyqlJl5NwO0GHDxem3g7bpbUMwj4DMqs9spP3P44KG/x0sgNDBBAEEMe2cC6I/Mx//v
Qc2wZbXaM7UhdSpm37Jg087tpQ8CzE3vdoPtR9+IfY9cIkRLSE+fOwMzqlsdN24TZ955N1ciWeo1
w0r25n2kJWsL5vJyjmS4GSWWedUnExVFWpWkEuodAMfmCJSJCRgD44wsvbPxo+0Uln9jSgayWRMM
P44OSsGYGjQ1Q2xNLde8vWbJhFj2YwF4BZd1fd9Q0AdnBe9fZXETORSCrhYwvsqKbAG2ipTtevno
C+2FArSPRYkpGcPzCzw3hfGbUQiiW1SAdJoURBNLrd0OBrFAkVduyhzmSXZ45BAOtyLi4T6a/+0G
jmA5hAUxlB9WsbQtGSKONMM2Z4RcMfklyZCnGnoeGaP19c5c1iFxz5gIOCx/cotv64RsFcIzDgSP
G9oDKplG4QkN8ETzYRStegELq/mM3XrWZLVHw8VUdRSkpW+G/0npR0ON8pDak8eaOGf512lF64CR
DNjW+GbnSm73X16Ag4Y6CVFYGGsMtuTy8OZWZgEKTPZtr+c2f+Ry7dGc1tVclNTeiBoOq8fJ8k88
hj16EyrCvrT5wtZUF10zKgY83Js08UFO06Z+SC6KTvD6on/KF3CIt1fzvbDKcfCuXHO/HOMkDXPi
zQhaHUnj+tAox9q4rnJyngHqAnABu0F7vlLcJ70L6P3r6pwycqpbghg7pTUuM/XhD2lDku/G4bdG
mVVwczXboWNa7/rPzu/2kUX+u6647cnO4zejoZzkZQ43fw1+LtYCUIOFbmhBYlV3mjGS+609FhYH
vcF03gkqbo4sMkr73LGR+t7/j4vIG0ATdB6n8IpY2TW4DDLyvuV8C/mwmzcLEvW4F/bEjGesqwTv
5Ud/+dAxdSLaS1MuazlTS0Lhc8xG+VESkYlu+71sZktCgecVrYkmsI3VzJmnSQx+75oRDXIch4et
2YeoJgn4ZIX/J373IbmWJgvZfcO1wn8ObO4Y04gmQNBqgF4mMV7k8f6gpuRAt+iZp8kh8x9FiAwW
RXYDN0Er4i9VdWkRGVf7xfCxIwZ8SzyP9crwj/lt/Sv1wE3n/1DOSyYJ891yHaGpfc9erU1Y0S7E
28ZjlkY1KgctQa8sTJArkbwMPM2ViyU4votM07/5SbV2lQSNo+SH/qMhD52T/cUnZCnSt65i/zNa
Z7ZhfYrKbvpV8lFQZET2D1OCFLVAgN8u06fosFaWXZZw0sK6SkP4eCHSt/WzTkxAJhGawNxDiriA
MuUCdtsDBsihgNHm0fXbKWursmL4xmfu4uzv+1nHEM1Hq7lQfBD+6w/ps4uG7eIp+/A9HZmWIwCJ
6WSdZ9YnE6NmWNQpd1pJUcdvQcy2b4t+E9MEYfzMchcFHObPWpxvLw5Qpp53KXIdI2ielRGsd8VZ
GNMA41fWjl/plTJMB+0NEwCgsfHsoKszEWrsR69S/6+5MwmQovukkqzjII0W2y03Xb+sxaR5sU6M
5il7EHsfjVm2vqWTJ9r1vMANpXVOUA/qiETzK2Lasz6LZV/1vJ/0DlCGnBOGYk68wjlFfaffV5I3
DErK30NH/rcanufYtkMYf8hlXKI7K7LF35wPkShklBDpTP6UlFFWb/Hs3VSyLiakwob2W3be258c
7S1htIWHrTG9ITc8o6KTIuZyLK1OYMEXtVJLP8m5pjHeUlYoaW88fePf/l3GaZIpgViazUZwkC2i
ekqgYrJPjcUc50vLrBb4R5leGYOFf1iqX5S84nV9EdRAWYnPr3aVaa749hqM1ypNCebflhW6Vb18
25SwplSDDo73tK+daUvlnS4FDfz92d8+C1QYNo5J18T6aR8XWAgoruYj3JEVDQ9mH4n1uABz5loP
GLlkXCfz63E3TrUg6pF9XsxNwVfyAGx+SAeC5LqDRyYP+2q9RYN8rP6WMSYVVNUXSklB97daD355
Gp5CnacBXR8swZghFRMOegfY+DfGjLb7r+OH5COAG1QvbzXcvQO8lEFraMeoXasb03b7JWSfuLK8
ba1YuMgE03v0ocCOa42+jaZhqprOEiWuanFIqkCL7aW85Uw1AtZUYb4bIo0s0UYvHNPm4JbB+XKQ
TJAps4NYosn3teIXSm/uuXcU/bY71qpP829Vfk4gVctdK29b76Ki8K1Sc+w9fOvE4PD/TSl2Ifuv
eXtTQZ8bzdEQ01La7832QShZHiZQyI+GpnqBe3xva2ZkfG/A3heLaaVNkDkHIYr8LQkaqkLj7Aj8
A9SFtyScl1ZmPfaDbRDdJVjNr+ehoAhXZnfR5chjG/BULA3A3jDasqZucGKvzCiRWaYXqOjxIW25
/lUxzyNYnCvNs9ld47+8danXb2q2wXKs+fmHq7l/98jc4XAOnXoqxBerbB0UnF4s5LGpg5WDeTFE
lrwuKmd1XCVi7HQYH1NL6EuAQfsosLnrxGGszl6TLc2c+RL2HvKz/4WkP+j2b96GMmBYFYlvBHqd
b73FRKjomriaZ6+ZnB2QQGIsVDyqPh+7k2Fs2ExdUw50pWHqq2Z1znNE9rzw2Ur6VFDqdatRt1Ne
a8fgl54Jf5QfOT2+3OfRviait/E7yBUMgPn+v2azRxRMdYqbg5wYeLtKGHMNyhpXBWucpXa2cPwG
sTvqZ6dGHwskAGVb4gLwBgoaQuYe++OpD0xtlmax8QDofq7A0LcsWVCgauLzMuxpeKMeVbqT1pft
IHIrCp/Tqrnau/4mQQv+iG82tVrriMGGU+Sa+6oue0LCyD7p+9C3cf8KHXbuMERu3UtV/nRk37g8
/Q+8OMRGymhaMI64J0weP2YxdGOB+YkMbC7bJ16KZQBi4C5k4oTOyoN6CYHfr1HIqPbKekD0tKPi
IBI0AqpObinEYHGANztCCLQdqdIQxeJDHZQJlWcbsG7VAolFRgyJ21uC+pgDAvRTJp7B7QOmEtf1
1/wgZtwlVjGVlqTpaHb3tTfU53Y8QiLXwDKOzp+pnXDk0vpk0Y0RAKCiSTc+uIlzQzg5poJ2MCqd
AKBT38hTFHohYrvUDcUnkzxwb4yylvbhlXYQcJd8+7qw1jl02rXs/LPZ4oad+9TYR/BzG6wKa8hP
3NqWzM0S/DgOk3+fvtDXlHOlV2Qblg9Y/JGR2w/QCcMuC1+Sf7oMh57VgPTDBytokD2ALpSG6w7i
z4+AlQTxc1BbKsp3e61QVbZZQT23M9zc7511zn/RsJu9OaOXoc53dBkEcrM3KWwGmZpoVBiSTumT
T4lBt7lwZgixJtVuWrqgFYcHLUCN/aIXxkTkt/dwOuC7G36gCMIGmg2yWCXuVyBbWufvaUxhYA2i
2Cz5K3o1PxQ6UxFVI/56vLuiNUOYNWfFowXeDQv0dcVkSGGUYz9z+kVPF2epmcs5Rmg+bIG7RNHN
RH2CQ149tCm66OBfnhl1gUnhnNNpVjEoQgYjsupn+x2Ycua070L3q5+xUGa3715H2HpOmuvbZriD
0l7ALq0fL+ixxDMMUY1mqb7UuPJu0H+3XTrX1HKVhNd9JlbDU3LXj3lIHQUhpLN9ECaHDaUoe8SK
IK8Gr3lG8oIi6UsQ8qjm5dZGpiQBc35jtvgKZXLPK2h+pkBlcWmdWgdISlfsBYsVU0Siju8DE/0z
gVwW9X9G9HFARffsL5y1FP1XdCnKNsukD088oTomMgaJPzcdFWeL8dbAU9Bi9ODh2t8eCctMeK5Z
1B7FGJA6y7W26oC+0Ym+A+TUgwt1yofXAD85RW4b3jDf42KSnDa9BmbnZwcSFXVCblvCGr05TmQc
j2qHVspfDv95Rnf5Ov+u+phKA0SAhoUnkKo9dQe6KwXtkK6tdTGzkk4s6Mz5AhBn5Qx9JNYMtVzK
VNsE/VfYESzmBZFr0jNUIwCSE4rw/crEFtdS+DzplpLuOn2M87yJQx0726uWa0voH4gvqXbcKpQy
a/oh+TGiD6ncP9APD7LMbXvtlctsRpRqHK08+gncQLl09HihCxgBWRIymhj3waAZYZ1TWSaHz7E4
/cCuBCRV6ItDb+KgyKp0GwPpuRTgWnmKh7/7hNeO1NqciMMWCKCIPMg0RDf0IUPQk0kHl4N6+Ni7
U43Lj6C+3DGzY/hpbX4IBqcNoa6PVffb25wabtrOGIq5Lg4s+A/d38xvagTPyo4ilv+LTP1OKMp4
K957kipT0WcxDCmgGslwEOauGNC/gBCflRQyaXmoNDOHSneZpjHlZviiNYwTTH/Yxn2HkiNyQL6a
oe0y+S/cR+edXBp5NiKUXqVL++K9gLm8q2fq5PikFGURkSvTZE74r2YA4wvTZwLzjm1kh/3Z6gPi
HbyfZee6Qt7eqd7SKgtu01BRaarWyrzfScYR0LtcmGM3sq0GBhRHxg+9uigWxcW+OYg44WqYi6rH
/zHUkGNRNcibDAs5luNocKLVUbrO0Fsl2NM4clo5howSIkNjfdks7heQboDTBdPGUo8V3zu6Y11H
L3sUBRYeLyckol2nREkxXJsrqKWWdl4sXtTNa+Ap0zPiZn0HYbKfllbFz5pkoUExriPsI+q8LPnL
y/GihGM5PTXP48hERKNL3PyedH7vuuqJyKR9RA8bcSt7RiN2LcmGAaVzFq+SEOHJ/b1L9EVA2bs2
8eyqSm9Sk8qQJYJ9+PrT5/RYrddWdEONEriywrAQ+SIthmumuMjDhP+Y8OKxS77xjofPhGEBvmy6
Qa296vzMC0a2bs3Z1V6AiSglWl4vseWFDDNrbAJ00ffsayPW+JGX2pjWtSQYNyWZIvviSXp5TRmp
LehgicY2t7Vpw36pZX+2ANS6d3ahXbOFW1AQq/wlWeYBCBSqKyq997AoQzRG3KUcKEw2ZmloS9Yq
gCp12yN4lGhFWWiJV54fd1PTftJGjDXaT2hFnLEiNxRZF+/HhuVQInFHPAEpm9EEzlvGn2TxrXBs
5IVSV7+15nbJY1Oh9+O3EHYAcE6w/ul7l7BW6CD2bwEgPScwWoaewExEV8yjnUpcMhI+XsYgEcES
xSiVT9vcVWE3eLTpWHwigyLIffIjXdzgMjNVjWmhQBrk2t1uokgpjlQpASK40B+QLtNaWoBNr0/z
HqX/oow8rYjtV9QfbG0CibnALCNytezz1hmxAMu4U2e4kk1t4wdMPtGE2zI82IaECL7Irq4GAtSB
EoHeB11M/tBkgxfmk9yLHBFj2Mim3vgXuh//0HkdKPVXGyyoeQpMEJSAULN60FW0e253NZUjcqSs
Zzm3AYJMLUT3sR3kL4OW2eNxfJBz1o5hwP4Vf7Dx9yc4q4gdvxpyLHED5/yga+xYBaZNWoIpUKqZ
tfFZi98jI2CL0mWOTLRzaAF80+SjqStrpv8SwWHFpV1rUhM2/zImg1FjmEWU5rQXCG65qO3vYcKE
K3I2/8OIKOU8NWyztfdU7YmqAMbqPcEE6rUKYDEVT5QWVTiGKTVcv7GjAsxJZpgZg9GJ+H/snQ+t
SjvMvw071LXrdLPOjBz0yCd+1KKmz1XznH7mwrzq9H091rOKd7C9QWYpB8e6siRs9FC1DOVoY/39
ptgNxsLxypddUfNC8MlcRcZLt4hGkxSsWEXRtf+wkARUXWXtII5qWZrrNwntOhz+p/pzgLJ7A0nG
xkU0fzA0NXQGmnGwN9ACJOUniu8NdW7l0DmILJe8k/AR+6g4iPwQcPt+x82NDsSP+5fHFz6nRzuk
TzCEzGQMzhKZzXHpeWCWwhr292VF/A5v3lP/OTQ783NDTHLf2rrGcE3wiBfbAR5VRSCFtVtMD+Hk
H4sIDzwrZhfVgijWxe00HOab4KrVjQctzXHd01TP6/rT7HPo3aLNZyTnc6XVxmaeci8gOSfbvGJK
fWW2bHjCJeRlPnMP35CFtQ8LTORwRrBWFpUJEp4AkLw4WgZmwYmBHSoHWaX9bywEtcbjYD2cy1p+
/Cf5cF88rOSq6XOkFB89ebLkeknpT1IHa0gOciiZREAGenOpde6mdV5yuMnn9NdN3nc+LYu42Lfi
NKMYp+g2zkqcMLoRaNXf1SJrCTnsViONKJuBJQYL0ML3Wq7yNIvjW67xz078aHPoQdYiDY0brQIf
lGsHwMdJCMKNNPSUKLCKMaQNBtHskX+ArH8Z823qFdPU2jq5ITnQA5RDm+4d2zVSP4qPM3KfkIt0
GAOM5SnviguHIbsOovyLpFcOQrtoyPNxbYryH0Q5mTi18nFsauQRQW936GsVsShrEOyqLRVA3lg/
1XtJSuwYeKtavIO2z0IMZnk8xyAQ3xrQaHC/iyUA1QKVE1LwWpYYasmXLNMQL3ZBB+ALaCXs5Uq9
UdMakOg6XKVXd6Nb750HtX1uRn75QVc1z4Foe96aiZa1RTDuMRl8ZTJTB1UH1hinP2xvMq/d4BXL
foW7KGjIoqL70EugWzphc1g3DzmJs621hByJCxvzj6qp89LIVag6CBSdpEJcywQhsy7dRDFfty+7
1dMD1APEnQlfokFxWYGAreLswRGBL4oPBYrG1R1IdG8UXG7R82/fwKJtVNbQgu3tgw+4xn045Duc
6uVVQ4QoKholtyBs0SRZmbRiWmnIfT2mAOaZYcW4kTDNeumgg2QKLLyjAeE9cT0S0AWEySOEjly9
sXNeNeq5Qx/cWL/ASbNltInTyMMjGV3Loem36reF+ZRGM4gzsjOtwSk9M41ImyNOxz9gIQSiYzJY
SJX3PssZFjm8vcErJmSekoB0MX09Fng13agAe0XrJYD5NgvI+7wkCpt+yWm0XV1Hoe5PFT1bQhWB
xaTRJ/xlykjzTzV/opCpnQdeYH5xiCALkV6drYU5ANLiAiLXGBiWoHQ3LvY2arTolsjb3eTL3eQw
AZQVGuEAPmaSeDTv4zC1lJsPtoGsCIoV2BO97QL+swyFV9bSqgX46F7KcpzTlmFumxSlJdyZs/ab
qjCh2OLy73Zxk6Y7OeBzaK/k2iRalreoEnv/FHbB9SCfaAhdHcdHLqkTqMO51S71nLffUpWuZ4/n
ZSDMKD9D1SDkeZFyI4tpisooMyqsJHj9E4RLX28W1JsQ+XF1juucne8pA3nr2wQAOAFDDf4Om0mR
mT7nui8+NjyuOYQSX3vbxSt6AXjBN+4ta8MbpLdLMbFCrk2RIGlP2cQez8LSkKQeBc+y5slCrH94
Z+7HT71lXl4lE6UbAqzNxC1BneZxTZ4cv8o5Gf+JRmNyaW71dQt3u442hcaLhBRI4aXEZB1ovjnt
fykjMAMpX3Ntc+80ZZqv3oStDrMYlD+hfgX34uWPC4QBhhvv4OatDDwgdsQjNUueWY7flzQNdbQ2
h3+qWlbHZYQ6Eg/X0IuDbbD8qbDWhJoU1iQbcakPxCE5KFuQFcwlhDOyTI2k1jy9NNNZaULdeySu
VSUyCHTvcd7EKRxgnhsHY+4k/dospxMvPBpE0TxDgAeVvfQllJDRiVG5TbGz/EQUjlFDT/LEzf2v
md2PkkcSq0+BB5WR6zCZlxAUS9OQDpo9h/SMn8E6q/0dS/iy/dSWaI7GdCVLzPBcM4X38V/QQlFP
2Y8WWi+Zdk2imAPYeyHHjqcab8XHPKF+bNhzL4u0H0+JnXysZcfZ8kEOyvreJfO2mVh++vsOw0Dd
eUP5ht3IOa7OVu9T9S1NA1Gg3J4CwivXg13Msyg/XBydvH7zYtRdBNkqB2WsJOdj+HpXJEPWAHA5
oMnWjqejgreKRQ+me2tfNE3rD9U1102w3v5u8CzEKkbgSWktkDGK9Ns4Afn07b8Yr80wQfBIcny0
izvvfjR8qGckiEHAJBV0GuzEllL+bvtN4jBUfHzAFQF8B55coGanjD73lXGXuAi5jhXwjwINl+cP
P0fGjCjM5AlTFb72wnZKI8piAxRiDgxqAIOkjnWL2gGTJ5vnOBr/cwZhXlUh3UQL2I5EjavNHHhn
BOiV1NJU2bo+a+8iVE8WetE4LHH3q38pocLTWv4+K7giAmdnG/lCaLOauvNannzZPS3XP2TvfnfC
16kppsd0O182qvMMrqpQURL44IJmU/iCzCS5mUh0WKgEVJvKiMFkNv/3Og9hmKs6/9+soeMVY9ym
K7Ik2V1HWDHXKdG0hnpsO6Z7q+8lWItKioYkGZTF/A6RHpIjL4qWuZwMQb7Dm36TlTwUR3DLxNjd
wsZYsLoJ9X5fPABgMALi8dLDcmM5z1S2HZCND+SRXGr7B8lTDfQmHleSqfhszuF9Xyx4gAAvipW8
lfOiGKaNyTDsYSdTdGV1aVvlZ9zWufSSV2H1JG+Zcp7lFw3ahifEXi1lBPrJ5gMSKxn1kAUVesOG
nzodHdWK2RrvUbCFCnDVU8oMezIW1kIQEFIur7vnYWEAOIo+okDTbEYujRHGzZxAwMgqhWiTjLpA
aShPviZ/3nTGPZirNcarT2KmXweLJrD0ro5ZR2oyd5eSDdsO5DZjVHRkjS36cF5o4hQ6Y8Dsg8jt
qJUo3DQyrlB0QpZKx4VSqfAX4AyHmbBPj/BBrRFOHvyiGRyuXLpRSee49E5P5i+xnvlISROJqdn+
fBYwHUgF3RQAFUHkQhCehnPSuGsU1EZTwsayOgLLAXkejvZJAFzXEdAx+2Lu/5DNY2ZIdCtUAnjm
xE92syrbKtAfiOTloiHXgSHnl1+/W+tNZZcE47ZfN0g04Dsx0YqXIRDgrc2C/LPkwgaz05tsXeWK
gjfwYY1kKp5/Q/RtU5+P5xxUwJksRMZdX6n/OFX0o7eRMSOr7E3+8SSb8DH8oBK8USXhmhc1p0RS
7I1vfWgAP8IdhrffWOODFnC/iafX/mlB0MH6vjOeJnd6gA7SDFYSAAx2u63JlY4wPX2bbxT5fMSI
+4o8zFuAqFr6Kdmh6N1orN58K/7hAKXGEIyUPKJPSmOqHIxpnzKtjDmxTH9VzVeBT0EnWIPkQM7G
spU/B0da0MBF/WN/5ppbvfoUmWq/qzHQEjFXKP+jEM8Mn5PL4xgVR+Gig1PXXru1plI8oI2LBuRt
DhFgYlHxz6YzfaqqL1GOHPV3SombBkLrT+qXvN7YKmdsiQqkDEP7Xug/DOKIyi8ej6RxF6iEOVhG
HJ7rOlTfe++ANjUelZnTUIPbauc+GQzxwVqoHQCCmUTdJTu/3+XgzkpiDdcND4xebt2qwM5i8tXP
UtVzMUfF//miI6EhXegloBk5dBrnaHuOlteIKx4sHAkzPCGz395+VPfvh3tT8GiA+8UX9tNUmI5z
wfhEXZg3897UmlJ9bGcIQB3GIZyljpXKhh4RqcYnxZN8b+IazD4T7PlbB5WTT8rzZiQmZtfGDyjt
/JVcSqXTWS6JmMdQWStM2O97GJVtxdcXlq9yo02+aODIQNikt+4CJB4IQnqAC33U6kdDiKpZ+hcW
x4YFLdBAPBjbiFT0xrhESwD7EicfLXY+L4l9Xnb+tH91MAgIPqGSBU09qGMFY9FE0eey3VxaKaIi
R3t7IMEGqyEEkT+nLNrHK98WpE5f00u927SpPQCWPwVB20kj1SAtCBuUXBBg7FiTnqduJvXQRH7v
Q+rirc/rh5c/fIeVpwQabLOExKxXoCUep0dysC5XDtT+QcHXbCSkMcDWvL5aoopR6A0NYZhrhkDm
2/HadTeHiBYK3yNNeJTbG8SR/OopOM/bUwhIDjK63HWU1g6S4PFLKswJS7j7f/o54yyI43vQXWk5
mRv7BQsdahuenmM/R1gzSE9s3CKJluZW7WvI2P+F+sOgESgob1zF4mlCk1tkFOYGxPC7exBDHbGj
x4S12kEHVHfBxA2rrDUjaXhflC4+lbUrehySYP0QrLS4QWsoY0bsC8uYrFDje3m/xPv4kQhDIbOA
s7ai+j24OuUQP6U4UZ6UnjYKdPiJupSJbaLO8QvtspjpyIBBrGJhaCxiBSs4P8BoqggQc8ZtTFgx
E8YuEkStv6UA04ymWw0MWW6+W0BfM2xQwkoY/o5AlZ5X9P/+0ZH0u0yaNRUNRMUDoO1TkGzr73cV
qn0oZd5HtnCkZHj+Aotvq36cRRq/Z/eiVV/egTS/GCAEehIqv3W70KSxjCNgMyz78s14O9yJXZkq
9wUhLYsevsrMR4A2vIdr+pngW/0cJCZA4zvUkQ8R0hmJCIenFNp1TdPFTPvzBZQ3UPnxX/iWKTAq
FSxvTVcW5bAG+HqfxsuuIkBm1cKEt9782G9810LAkLcQQDv2ey5mZW88UuzunIhHuC17Cn/YJEu/
6Z6WQvPBRY/5WJ4U9pFY4vX70vo80ePatoVfh5bGhNhN5xzgP1nTNrLYwTMjIjUiEFE20oXv4kyE
jHYYtVvWRo0kdJAmuyZu/bj6miS5CD7PEATe/mO67fPX8m7AVGZkFdwmIe8pJSg/vL+zbgMklrSq
K6324qcD6IrpxBI9/2DeTPSqK/sOcE65TdQHDP5tDkMYjnRhS584MA4aH1JT4W7iq+We5Cwd+WWX
BcbLOU9hX0sJZX9a0rHjBZqkTbj9Y1qZsrP7opdiL/ARi2osL/+I30YpnCNO2vgTn32TaoFeN8Gk
eveuF2MZrM9ymJ65FW4ykl7h0ZThqKYZSqbIf/eRE+j1uxBqCsBC4iim+RCZ/SizVD8lAr0C6zr2
0TVyUrJoM61j4eu4ay++MLuc9Do/uj1YjRxi2/SUOgHiwlT38t+nNz56phD8elW2Mpx05T1UggfP
Rx0X00bYox35qAb4QIDf5V2NvfJhBO8ap5kTcJyTm5oZv3CVT5/53jx5474clLX90W8NEB0jpsD+
ZBvnZE4ELfAJegbiWNYb37JuYBPLGawVjFcvmA2jxTEZHs4cu7oa0wYHRIzoMHHbOicEjDSJYVl3
qhBdeKu14IofbND3vKmRhVwCLNe9RKAgK6zce1XYZpCwpuU9otkPlhEILiVgGOsMQdBHEAhT+ReZ
MnY1zvL5f3FI0i09/yvF7j6rrflvz7STFx1z0WFSgAaTCsCfYlH3eC/v7TXd0mVT+ooAhAW3ti8t
r1XuiFjWiJHrygFOgrzNa6yPzsOC/gEgWR3S2gV8YtNAeQ/8tSkIC2xPtHw2WYS27230re8jYsg6
eWPtiPidmfSsUQGmZ294nTN2/lWd+tTMqky7ycURi7p6jWkLkg1bBM/bfPLjPQb1C0PjSKfC/NZx
3qRZVd4AD4X+8LGTcrzV0xdnqWkVFQt9r0BhKFlcBuo70Tl6cTneMPpGG/AtdbnRe/I1TWO90uac
62QaJN/enem2BEECaufoC7aaqfJu84xMWQrPLLFWs1UEFaGbiYt/+adRMBPlpy4a6nUYEJGMDqWL
rx08eiTUwaCUso5fShAZBkKv6ZUK6NfvVZ11XYGBG31Q+zUAq+4niDHVg0xd0u5D1H8pB2AW0WEP
PQ7MuY5oMFzNnV3v4QqXiLJ1eZPIaSKSVfPL3Vu/mHjeq59CGpxgwTMxfFU0OsnidTavRd5GrUiq
jAKD2ToWcti9HriVN0plqf8VHgrQlc0Y+r1diQKajgIHYWrSANEEL8TE40Y4bSn0pX0mSuwfSXtG
GNU5XNdAhXqljGwUpCHXAAmiM1e8t1ObANjucVumGoloZ7N0cQPNOweC4oR/5p+B2/RXWPBslTzM
pZoq4+7nP9PkOQPUbQsDu35HSzjQcZuKAJFZgBM8NEFv7GAF9F3yNBgpmgaI+iUFcEKclvKAuuEe
Z9BPoCwjKDoQdz8d91IOlVsYrdV3YTAIJoWEkNWGfb3ONwd5JJDUFbzvvrvxUTXezrMpZrHbZnUf
pSS/i10+9rrEhm8QZM+drLOhHtUDRS1xZYVBu8bhrU/eTIds+04wZdPunYlPXH0doIcbMh7BcmFO
Qv/7Y2MTlB4APqfJ/nYAT+1jXNihQDCOBrnkGe6WaDHDqGKTTvtWcOmNmc5hutsSJWJXN5K/0WzV
+bBOx2XoQPvX5LPLyDzFm3WuvD1LqAbC8qp7pZ2j94ij9S1Hz04eh7Q793qKR9CNkd/mlKgMt6bA
lAVgMdTMARhHSnwEvOmtEDru4mDnts3FE3oRM8zvwqRVVwiguSjz2ZgJ153E3m7f2+OVj1ZqsG6i
TNqIeL7hQ2YAr6387LanruSz9ui5DmE+q2pSZ1U4/MXJTHOOrXVSceuAPakXl1WtW3LihVuJdu9h
1J+c20NXQwmJzuwTSuLnf65by6IWYvaoLmI0u4jMo6DSPaMr3rGU8J0wAJW7nujX5RL7BJspa7XI
8uM+D1TuMZCMo2+IxJO4gtkR3NlyGHYtoSROET82uK3Ifg30r/0dWAn2VoGdKt/oVk3EDkuu6yl9
TL3TJ0QIAt2ZNgIg6fj7CCYg++juTSHkFQ24EvJv4vWuqmT6h6Rk9+xwcquALgg2pwl1+SoDFlIg
J8rfXEiGiAvlhvVYtKGVSAqX8Ic6J4ze4xrdHKumdwWphoQQMuIHg2s+idKjACPneiPCzjfQQDHO
CAMtukFexjXcQ1pjc8zpXk2DUzXRsmUbwcU71JeIoZrMVO8YSzoyUgyxH7kNZsMNu7ARCEocYWD/
gR77FqdlM88OyoysnupRsmvG2ljzYoNSerzP3/wNaKjr8pF+GqWZEPhfezwFG75LneuQAJVtsioG
tcULl0lGpQL8hTIOO30lQ6+KTOO2FkkUbx+8WTjTWK5ic/mc37okVx7BjHt3YdNU0Ss7TkLLYMir
uGIvCLB5uA2TFc+0hn5hN/IlSuJyQH5Izi4ov73CExyjwrSBuiaLGzH5bjbVyJR/AclHfHjOYIEn
t02jvJ7oYGN/ysWZTE7O7V882cW5dOaZy5cx60TuK/7o5ON+xGOmYR/lLmq1pdtLYnfbmrvctK+a
myPQlGbWSpLnWd2XQhx2esuxCVjbe6+gZFmwb5IoeqEJRT1DhYhI7Uv3ItIjVBoIGmUDUWARnRxV
1EWSZWwo7fb9LBJIHpd9NXPooBZrQ3XyJ9g3M42LfY7LGAcwFrfvuMP4Pg/ntH7yBSruyDfwLwDv
rYOmxoHlS9qAZIRZ2v/bYUFjdzma6mPL+M3k6g5y/vgOm1cfWTSutQasED5hslfYmKkucuZ+9/BW
M6wlncoD0FtbTu2AQQ8FU2woJIli8usN4XQCfMC+72koN14ay+XkFhKGEuYu9GrUiMp5AmTWOh4g
mC0ruNjdD6iuL/IcvjZ1p8kw7UAhyLhp66jr9cgmOh60lxZQ9rUM88iGO95ybSzev3vb2i9YOSfe
tHCL1XXy4h+Fw+s/r4jS+AWBFvWTK/H4Nv+9ReQGIRf5cTmsinSnypxIVmPX5msG9U+HRwvpnVDG
s6sZ/r/+cmXozLreF9JvhqQgmuRo5I5sYuBTKIMMFq55Fwn45UJ+xJqqQK+QVtWdl0PeVSIE9vzK
7qCSEdUdFJeMlcW4IPXcjUh6U9XwXWUVgVa1fGVYx29DMbOmTVrLfjwm4mIYj+T5h5VkawWZwH8n
UVuFAt/X4WOzjiBmlpC/QYsuJOFWWKxkU88ex59rQICjPPKp/8wYMPLEGfO7/ZAnzFO0HKr203c+
S0qjbQ3r5RGF7B1VpuoeUG64QhmPEhjISJ7UaQ+usRr3tN9J2s3tTOz34tmKXcHOVg4VvwhSX1Jw
YEvzYa/+h2JfvlMPL4dZt7kT+wpeuI3ha8rx1rFB0pfL/Mt5gnaFlQNbOXSFGBFKpJpYbyvhqKS5
tiy+yLw8XCZ7kfv35f3h0EZkjnHc+srpOj4J+kIuQhYkDeNyl1oX3aGXr0fpZXPVfMqZXe05lmlj
B7/Od6729mFuKXpc6RRiPgC/OBJmIxeMWb9lNgeBthCdco+ZIiJ4cPsRmVJJOyDBHIMIm7Ub+Tos
4JXr+ZXheYXzlsl8gogLdsY3U847kiowgFcXLfw0PMBNw+dCYlqd2dG1OtJzITmxMcDs+pdXYQpA
uU1t1sqswqcN1lr2HKmc1S2rH7PJ+KECkXma7I7aRqsLhq0uy5ph6ep7vV+Z8WOhjwSDvcASueGg
RTxx+iPt9fhtTSDMySa+KXOG67DxZ/gmmif5ifRJzv0UuP6FZI9CGpRDLO7ThPSAVNBXzQlW2bHb
5rWw5GI3ROhNb0sNoxj8fZSD6CUz0MOtVQU6F3+nARi/4Abp+YvU0aYZD7cF5EbKjyfTc5zr3QWV
DqtvQ2Jw43hyVceL3R+hUdfxRSNl43zt3RLjHj6pogoSOMePxMgQ+i2AS0hlexIaoE0VPYWuUNHH
povkYpS7Gt7td/RmS3kBvedRIh5DL+ZRgciMbEIdlizbtdcYNbwBeMP8wA0Mnkp0KO35qZEwQRUF
GVNbnL2fySlzaA7M9/Xuu5j7kzC6hElRnNFZRvSY6l5c0H/yXPltcn6udQk3QOP3bE+/mEBAuCvl
GYqvFF6ILWBBwD7eDriCbU0TajJAFUu/TnXSQRD/ltvyOySNImJva0sbAQfGmlbzx2Bphz+2Gn3w
AwP7MFYiY09N5IengBhppQXYoHDtumgK97Mk07uXJ8T/LMT+ds0/rrjdeozeT8iQZitSJeeBUtW6
ZaP/bUrOyq+zbZlD9025ZEkBzIVIkARG/7i4IL0XFY0JKza3yZppYK1cglF8/HCWIk/QjLn0qoax
n7kUrvoxRZ4oAjwOhMkFBo4SGUYqo/QcwF+2BokqNpoeicrsz4bm2itiFHQOBEo9QGWe6THgU/Uw
dDfzYx4IZhdNxMuzciXShcqeIhJM7wRumWA8hCowHkPwICAcDmeSm78gmoOegzRzQ/5C+1OuhLCF
SdQ2kHBj+bt01rg9saZ6hmWjX4zBjab9NHeI+0cRnanpuC6KTf6rJARiGXV8SVmNAUuEmiACxMuW
JuBTFtfiE+90eB4y4QS1pEtXCHShD4e0KVerBnYblCdLha2niNX+ftk9DmRmwn/ZZDwWruCilEVG
d+CnkVQy5sQS191dh1aOH+Pxv9kfHvzz6w6bxR6xKDRk9EB+zMrVsxs9DbkcToBwEtb/zz24tOOa
dYH0y+6bT/PXJsXh6btYGx5kSyfoTLjXnReZc5DFKTfhBD2aE5+kA2nguGxNpaaPmhSgO8rF9yNi
v9L3IArkvpfAcrMObCzfl9kwgKbg7bL3vyh+TyU3bKvl/EqiCfJwOLwyT5xAJvc+LxIbxO9i9/rX
pfI6gzPTziYDXFbND9otMYiA2toaaMMMR8froXUTFzY/eIxM87rdOFOV6Y2bym6fHZ6FQr574att
HCl9U6WAQVVN8BP0HnSMqXrBkgiqKeEOQJey6AP21M5YWJILl7ZYISTgoiw9eDQxSOBYQmUp9ahQ
rj372/QXZd6Urmgh/TZfdb6vVnfYNofUuAqq5mne8LpUB9e+VZWt7jsCR03+eW9ptbhE6uO3Ecp8
/jRKY0Xqe+d9lSlABvFmssTFx5UCEZc2i8RiRxF2onUmfNJCHsmfpCtKzZ0I6d4z93DN7x6g06Gd
Ai0HvBje/ws7KAWT5BlKxgGDZty3BxpNlhF5w/iw1fh6DlqCi4nV6BNvTgwtSZMwjgoQS6oY8jP4
gN+FAmzwagNyIwO7AC5pGiRlPOR3khzqXsSstjgHLH8THyKn8vOqanLMDsY2nKsFSp5QIR53kzan
iemoaTuJeu+GKx41ar6qt6EVZsnunHagoeAUfJyd64DQBVpiRp+bpe/7kxEiFnipaShXps0qK9bT
Y57VFysy4mATV1NIvnYGlwtowPdOd+TFjkugwVdwzk6j12wL69Fs1VomXHlTZqeEp6oExNQz+4/v
Ww3JB6jBasWPaLJjnuaq8cN3T9g37UFlhQ6l3ZFLdTDmT7jM6HuPLylWUciESeB0LKKOLrKWZwU7
iDJ3PKa52BZcRJ8ykMEGoR2JjAS/4iFe912lJ5StH6n1sAlrkWpqtxk7jXWKQxQ42/lISoiNZmva
Ny5GP8WIiJhbOeMVBK8MLWG3mojdak1jzuPHe0imNcd8qjxIKdJvtwyTYyoH89etTN1Zw56HCeZl
QWBZ3EuLgSL/b6NXzTs/oX9ZE84zIYq8m8ZcUA4gJt/ek1yRMG9D8yZe8EvjLZMaBV6wNnoWEPf+
bde8yW8eovJ0JxU38K/r8TRApE2yN0/2NVi7WyZScbowQ4gX83cQDc2a2FPVzMwOH2txY0I+FY6d
MWOoudE5ZxP+PqsgMkaHXV6m5SRZE1Jb6pOkX3Tc6CVJiUg6+6LpAWJIW18RiimtPZCcZ9ci41Dz
yTI3gq85J1LUbhleOMf0+AvR97mSm4nuSy+QshgjJh/gfvTQhEmA/ip8MNUB3QOVupNJQp5QIXsf
HDSgknnJX25s/oCNQnwdYMD3vuR+5/LFASdgblziwhrcyzEEIPTE8/z++CgkFPGwC13/La1nW9Go
H7idrMda/6mX+bPVS5wL8YhxyB4J8Yr/iVBFNw/EZesFPwINqhbDJq5CUz4IdKm7CBEKUeppCef1
hnuMznuHfQ499U0IFu4aOs2IQBPzgU/iqsyj6sIvd8Av8rxJ90Me2xNiiStYShS2SZ/Xx8q5qdM1
HDws/HSbjASvFQSXHLzU6ccmGS7CY+1/gjTHxexySjoeDet9l7bgeoZA86looMZ632/0RL/J2l4U
cRjFimQSCxUZJDODv4xOQFKpnKD02SY+VkpwvOvYu/6NTvBLtZKVbPU8pATqmJ8Y8P076+UCRxIx
v6FVzkDsSKTM9wY2dAgrwZOxk40/GusNuyFChlBUb+/BiMongv/5SMGHD9Y3+361BCZYebKDA+TI
H1ki+YqpHFSO/P+pDJGO0fOVnR5YsiqDfTIDxfw1C1A0FKIeSctSiLhwBj8IQresVjeCGBQU45vI
0nG8/0AgcRFhXaMVaoikVOHWA1tqgBL59lTapL3MljvjzjpJuHUxCTCTt1kDBOyENneNd4jLeaPf
Yx+80gaZywxS6dznL9Sw9AzQGwdbh0vsBv1fhnUym8IwwZNQPhn8Z2ChoS4sG+uCSfpG12pVADuW
seQJQCTfxz6AJbxIxmWbK+zboRd1fKWoMvPB+9HNYHKPhncwuE9Ib70fQZd+AynDhWDZMbGfC9n9
za+rsFtSX1m8lfirmy9r/GcU/KtZ04LpOZv0cHx4gEWoaCICxV6K4bIRnpkvPAczSdwYPUXnqjJ5
smh7SWB4TRZ5HOcpWn7+vCaAknxpStkio8aAmuiMWlMKd1BfsPOjoTTkimFJgmYDhkBi6axf2mx8
N9RHxukIH+JmidYY2PLrGQL+E4un561pwhViGLvOQ8S8l09YBuw/SIDkS+2XutmeTpgAgjPiYBdq
gbM8L+f2K5NYi2YVyBTn3iwMPtwTecuL/kKktgGJtYviys1VDGNLGfsQnLXKXCxEmI3i9G9dC0Az
A0z8EUDcVTbjHkMHK7p8QaHQwIhOj5gLzuU5PHSM/zY9wThSLy/PfQe7lxciA8r0E3uh1gQJVKc9
rg48WdvFhI31bKxUeFD4sM1C44SulhNBYTbn8iiKPJAMhMEZ8rY1qqoLXBXl2TQ3LhVuBjgtnaHU
FUEMepxvwgDUXXCxEfLV9DqBOmc7xAvV9iVYFJI6AJHh3UKBK+W0FNuVdv0HNFTBYUroadGHpulG
w5dHIaR37wASbQC5DhdtC729On5uvyWjBtU2wLJ1JV6/gjq9u7wk6jkTxK+Kkr+QUz/H3ADKxJ6T
PRyttN2tJUSK0kQbKbf4TZqNJ5NIwphswlFbXKQOH0c5/JRK9E+WhdLWWZukfwARS8lOzgva3V7R
nEWo7/+nNEq342TvqiF6UKEfaZkPdXjMiDtuxSElT6aVM/0RotJDA2ro772SRPcH3HeBgHHXnN73
Aq0Aa5XIrl4FvdpnLfwRg1X5++b0zZXGjC3hstIcWn2JmIhMzwc1lSOtC23U6sM97sWy/3cpxi0c
zjlzrugdGpF0LhWlvz9nOqL2ssvW5gmz9uXorKQ5I0g9YIoiYDh6fWCnQIO9tP5jDFLfQeP577tF
zpuYu4ZgXQJix6pOXFVxmIqzMXJzZhdmzMnNSUMtk4Uw3OO3Rwj0G7G1DMAuGG/dCKrozxXYivZj
7wgdImDbb0MXlPfTsYFfpXp8tzFqh72cxSzbNJ37Xtpd5whXZTq+n4nFK3QWDR4BbDyC0KNlIPBZ
8TXAjns5T8DvS8cMcHgxWmh0wp+DGz+C52x0L+glA7Z0L3kJCVPlnTE1QTYLBh8llhNDwPzdwlgz
ed1BPwnMU7gjWFk2eqlc6NPC3cKlcIwYEESDCPXtl3/gaH4+Y0boyLXdgS60MbBb//AzluWgB+ji
Hqr8P8C55U6yKep5LfY3yIH20bgX/zkR0MWPuVjfk2y22VpKJFzyHAmnIUH5Mrp7nzMGiemV2Jc0
alVO4qSbaQ6i17oJoprfBfq/LZtmkfAAdkB8d8JWEmeHWrCkodsaH52K/LabC/7BZdr7KU0b/oyB
AI945C7b9/Erbgb6E+MOgrHXNo/YOnQhYsrWJxQUondWZgH+yVP/8/HUrPWl0NByvEHf4YtdJegq
lbpuacNH1lbj7Ej4SV4gYvLu8ZcmryHpes2sNdw8LOL8GyFXStcn+mx3E53/m66b0Yp1BTOWB4/U
MEe6mcQmXg2vF3VXrowHNLq2Zfqjloe3a+x6R64Tlc15/TgBZY0RGLjO5WI1xPDTwRbD0a9Lsmkr
BDP9auAxHeDsWjwFpWtj9QKc9PuT3jqHVQRC0HFvX5rDf561k8cV7G501MTajSk2zQj3vjMrDgM6
6Gy3wuWJwWZm2R3NP6o9pWgO2YPtZv04zge0ZLuFvHXHfCQpbS0mnqpTzwOWp40AC+pQVSCDx+Bo
Ei24NmtP3hudOiZqntf0WiZnBuZSw2YQfLgEw7J0bVurNSrg0UB5IJhRDk4YmT30ULDNnC/S0dtY
zvTyP3qsUX5PNYrDSZdArkANYyHQAtlOef2uzR6432X4fItFaPFgf4NbKHCniB+rJMf9mZMA51sS
NLegSVIFxfuJgIROW9vm6xha5hM3QUmbyl0RU2GJfJIfSQvZ9Q09l2yKsbvP7EfOIHRGuk/tL0Lt
F30vQezFoErBv1WPAYTzFn+IRLP64cQNhSMRfxAcmOsC9skaY4L4wbWF66GSsW9RQelXV5On7Poy
JaVgS/z51ZX0RZ7VaPvEXeQtM/GZtiUHb0fgBuMUTFzxPNekJbYhGicEtXyVsLfT+kAduh4ZFq7f
A4mga/hBMTcXmI2TzbwLxcyua/lgyPlBoxOinEjQu9eyTJX0bhuaHFUeHVYV3103hbPBhj7CZ0eU
VjCImMdD6NuGN/3paGX4WUjRw0F573oN0FLXbS+RD0BxNlSMHGvaSYPXSHIFTlPVRbT1BrNUnMGe
6O4vzPMb491fxyQ53dA7FB6uo5re2RRZ0OPwQjPMAVIOerdKDoKmMusrxo/SSB18u2pm24cY2dIw
NagVtFUXmTNNcbNLZlKric1jTzcNFgdUA3A0zvKMoripBJ1iOaRoQG4wFVkZD+4QPMrPuDIo8pXX
O5TjxTsHqK72CNkZiZ+Mw0o+IDvlDCtg4heHFdBCJrF1MZ+K2Y21JwXFmrHFlTGlRExr2TvvcEFl
qux6fV0DBebTLO6v7aMO3t8i9kkFua5Fczwm/R/7vmjaX7278YDr/hdjqsauzZDwFmB/Wo8Dg7dA
4rocKuS7BDS8acwdDJGDhJBpTVRAnyP63wXbEhap5uytoU6JzhWb7to+IYRw3oNdDd+Lhq9t6z8I
hSIO3jB24rLc5VtJxlhtdOKXNX5CvoCLHLIE7r15wSo2YpgTGTts2hSpkhBr8R5NvEB4Uw74JSVW
yQ/KMV9xaeWCUL6+Sm6cHgQqu0quNmwdfvP1pRRX7DGYFyxihzXHllZMV63V8EcdxO8lcPmMB5gt
4Eiw+b5zpy1h4QUONEUpirzlDfAxY4fdPN3HpeYJLQY+powQT5NXlLX/j99VqahRRIEpYWknXnoa
/xaehrc/ig55E/Y4uub9Q9J0dop7L/VBqNrLx/gvi5FUxyNBPFJJm92DdKW16QXtnscP705fAWe1
Pqq/kzTIEo8oTpVmgurCrqygTvoAHsNMjV0+VVzfys+nHlTHFBQD8pE9+sODFv/Di9aFM0x4cyky
aLU3LZl7VgEKimaKSJHbaEWs+GWDwn1CSbQ1gn0mh6/5Xsldf8yPDx66eMdFHLmg7o0/knB6854z
QMNqXs+P9WqMEKAUiX404cVCVepkDD9zzDp6ue7yoX4s6NVOHtxxk9VGPaAuIPeIYwkZepK9ey05
YvuAOGFswhyQYNnGc1acOPLRSzWxKjrstTt2puVrLOF3yRYZe6vz4pJYVFKdkQs09JQUuKqu+NXq
RmTqgwB1Pqs+RlFT487mRvOP9iplqNPNib6xmoN5M40wTzcDW2Bebti6HzyHG6Ho2jGYdnnogECT
Tfab5TG1i9MWS5bz8FM72Jl0fHlzQySfosj5QdvYRK2M/FQ7t4JKbbE1+9MArWqVth+UkMrbNpL8
9pcGGT7+cfWlDLrmp2A2R1j90p4E4b7CajsRcv89otu+aQ4izwE263WymMF7a461cEJDRtXVr6lr
oiPBUp8t0pYaYFsmz02tUoT5QMbx2PGwjYF9zkMDyRzrGy3IZYdQhbvbIbtGucJj+9xvoVNC/uJx
uTeRv0qKqiALhvHqe7BLNBnE0O7ybxg2TaLJVkhp1DvkfQiFO5fVTTpw4kUj2j9H8QxausCprpwO
LmmYcCZZicc21TOdB3kRb04aW1Bs13+6cua1m1x7gNqfPck47hSswHL+sLeqF4lrT2S86I7UeFEL
4LD00l1QV+PRrHA//RKnJr4pXB2ktIBmzQonL4E1xwaYkHhxgkL1dQ3T6tw5EENChxa10RHtbZSE
GspQi3rCU6RsmougLvXuhaOIJ4ha6aeGSN3VUzGqBy8GPDFpRf9Ayq8vl48nwrQSDgZbHA+71D9x
wqCtQkFeb4bO2kfnqS3qNy1XE3UuBhZdbOpkWHpgORHaZQpGgQRWfbJrtsjpcEnRt8rjGMwOlJka
+iRlRnQuOKVWP9QwnSrj0nXyqhPZ14iSJH9PL6e++xc7EZOlDvUATZPn9sFZJ1LAt72DKr0BTcjo
McdVsxrFYew2vrKoKF0wAW5+2o2DdhXfe7UF+g6es2UrIMyQC027y5ZQAbgWGCJA3Yo6JbIEuOzz
4aj/ZCl4fLyk6CBaqGvWA6+qz06s1Pac9qV89wYiTTPcPYedZOTan2E3gAF9w/a6ssAOlVYryRRk
qDMRJ9oDZtXaQBtgMN2s3joCMclCwq3J+XmDaaAo85XWZequqy18qGPjGcm3MI3JjrJm6s7+hGzk
BxxuQgjgI3tNfYzSMKUkiwUk1zme5ARYbQof6ZieqLsmRsZLtIpZHpu9aGfQH0j0RmK7hrC7t/7F
TAs1uX4R8zhi5HaTck8+4e0oFqPC6RNYqd/AzOVcye520G5IEwW7nQw1i2c9Pid33jMGWigin8tp
7tYWXVAT2kezSNO71ryPLJd9fy12WzMAGiAQz08AokxkKjkAMkvorr2wqu/tJlM8tlu1lYWnoOLn
L2sz1rqfawTC+8diCOlRhN2jCYdv5wpzpCwt7qKWusCq21jqUDYtPT+u1a+YizXwkXPruIAX58yQ
GhFKnLOz50BdisxjgbSMHLhk/lrY1imvf0jVZEaAu0uqyOWpTnccE5qWjrelb7d5HwUtT6biGjyY
G/TE+xzK0m9D4eI8NuEqiLBy2ENjOcPxt19r7SUVtfnuD0hDbZX3yFV1YMNCHiQl1KzcqDmKTthK
OkGtmEIaTMjmmmcKlCv8EapeCCcMGriZfoohQ4dOzVNM0AgGdwFMdG8h0Qsn7F+C6LivMIwOK3es
ulzWahHXU8IUEy5ijZX/3oZ93tgYBOUUN5yTQ2G8PY2qsJ11TCUcPeKOXWDRTieMO4k1dk1ehOLH
x6fXtO9/OjF2FNXfQG+lckdQkzLTtos6zENlzqP8NugbIjfOd+7HyYEaAxqMck8PM3YFkOPuldbl
7Np0Ywh0LEZ2x2TAHMypFr+bG6QKDU8CQRSh9aRLxPWLU8hyV2b2xVdfoPqKy8Y6geqKmxAqpLf7
PtfIPgeNoBsaipIuQIB+pHvviyqVMne1klSE/cDWUueq22E+wabQUZo/GWymQITcPu+IEcN/mvkI
IXfwX0ZSG4JqkdEXmWgSBmRKipEYIDOK97yv00fM42HFf19JduOMfi/HD8wbzDXb81t/lZ7QEwYY
VfqhB9N/8KT8jU4wBYyAdjq1L3kJDnFmyUVU3tUZLs0gLXB3/E359iCWz2w6Os+z2hQSrKgjntSW
UQhxdvmmXLJP0TYUtJAlgMqRcWmAka72Vcep9QfDNIEbeSxjl8X9PmAMcAVrh5TZw2FFZ0ohjFRD
AmEy7myIe6wGQxUyeKrCj7fau0zZlzajRaEi+2m6Ps/zpY8uF1j1aWQpH3d8zRI5QisvHmzHJU2i
/qtjXdoJRzpxX7jS4zcviXXiXzxbs9bhVYK2XbPYJaCLNKBSGK6z7BeNMtkI2yx7bX+tSluC0iM4
QSotscSg8Pzxks5f7WW0izsmO+n87EFVxbfx2s7C7D5mvF249BDwYTJwOoQAV/YiqFKSgzbLUyED
Cgvt+Py7LDaPm9DAyR1wf6cVdLBejncPtzyFSo7J1Ll1tXpHHLVDxcHOvt1BO0FiThWfTXwJfUhw
3mVCRNMMIplZTmD/sAXaU9j2QqIUfSu2DABhDDuvriL0tWGW+xRBtLqISKhbQDOZXj2lB/z8C4NL
CPTLnwGb64gTZw/1Dyc4KUrk+urz+NmUbEyIi8QL68aFGYqZxgTlkF9L0oTTNg/uh4BNuDvlIcxk
coDlCJILpRP8RfJ0JyFE9oNBYxE7KCBkAWU/JDSTCdaV13n1K5CroRkkhC9tnowFnumkUfK0QJap
7Yp7vwvYCwaWmKUvy1z7lBep/20cwvj0Eysi5E4ocMrLGhalERSJSqUk0pfq3F3qizpdr/lo7ifg
C4E1ZG5EQTimL8MrT0UVyerHbFGXsVDS5q1H6N+ToYPuYYWHydptwoj068iWCqmDjOBx2whhJwXT
pGAhZ7rm7RCxaqPT0PYfFS3ALrnFSDZRF4hX1pLLT3o81cRDI8fIeBg60GtsTjBxZpi4OfnQmEWm
XL3IBnOUAHmrekcoxOsrZ3Ato/AlMaT+82Sj1nwiEtAwNkpXy0bZF+5wr1vvaQBmD2h1AN08wR9m
hJDQ+uBJCEKGXqhWS/0+K3WXlKxm6r0dytjaZczOlNf5L2uwdKeb4IUmkMViKNBs1h13z8a53OdB
OqHqYp5W/ccwpY3wZfXEdGwEa7vfEUCv4jG5pi6bblFk1gIb2ZJW3z4ynz51CLgreu275fUWSanm
3AfGZojBDVNIPoaCpFFP1DtmLQdC89ftGv70aB14+x169ZoorXFhjlyKErPnZvZ8rooO2hHM05Cp
0VGDvynq7j431uBFlF6ylDV1PNfEe72dP1AFzd5Y1ALOFTbYaWBm4PZhJxBSQpFsDKZk4TSuzIdg
Z+CCOxOfXaF1AhF7WB7fjYH8gUBmRA9v0VwhtySKTEfH42a1hWpRCGqlvzw2eOTJW7lQNnxtwdgC
S9ydJZlP8lxzyNzriVB0n2Ofp7u1+ShAhHypLo3gEIcs79tM8TDdshNdna7+WdChOHkL9THOmARU
Oj4sGlmEFxxwn0IL3xWgINKdYD4RiO58quC8jy+DmvWeXTt3dhAaefSPlyd6fnhnc7diuEz6jxQR
ql6OugCZHRqcvsE20w3lUu4qiY3ZpUAIxIehq3j0a/kZAtRoD4DoynVFocIA0fivibpIqk9IhVtO
S2KDm0e0Mw4eeIC3x1pQ+Z9uEP3ssC+Rhi/6h/MyrP2snWoOo5H5I80iHNItcLDhNs+nQRlNKMk7
3q66S8meLCa/mI+0t4OdXkoXLYg8CJQ9PAv0q843cjctL81IBRXrQlfw6d1KBuCL88YN3J6ZTs1k
Mj2+Q4ST57lOFkFgJJ0uzLhLeXMr5MWibBP3wKDqpZC+7WO+uGYywUhT7ZGRItd6JjUUEAp52UUN
FYNGyOtv6wTXziR1l5cGlvyY/ua20ynyapn4/v7k8uxKV4xsYNVCYnCYGQRdKkW++gbFhrfmsNMG
diYKGMeEwspjoidG7dp+oSAJdxMI1ISsIMX78Y8RHarvcLGArBX02n12AZ97FMhxgw+JTvZ81Wlr
hVO4JfV9WW63R/cls73ao1AIQOYYOFbDCvFcUSAFZxD7y38pLVxOzGFM8wD4Y+UwRVyxtSkB9YzY
x3ML+FG7iOKP+YAlDdjkVNHMkgrKak4/O0OgfUI19oZKlxY/JZEYMaZXr4xoyuENDW9ERlxRoxUW
YhX6qD+c5m7NnvaFAKaRAUwqPzFHJ/pCr7ysLnGbyBXGqrxPyj/nSjys6SYvEclzxlPfCvta153g
v26SLzZLsKuvZp2X6AR5m9nIuiYwd4+rN0phyfT/CrBuV6EhtvHOR7S+DkTtIJNQmDpon9t2K4JZ
bD6KMLTSmM/A+6uMsfhyfoB0BBHsfHAt01v0KvbfRHzNoXate+xq14hoYLBQ06BRHjBGx/8EYzmj
MNsEO+AAsmYUgd+xzCLh/iM9sHxuh7exXZQQCrTXCphUFnVchQXtpotvllwRfO7ByFJ8qJ8QNq18
+1FbZClcWNJ1Q/tBl7XIU0bUcj0YQJm6z1DTTFw1EMx3xexEALW5UHcbre0TpsYHHhJa/Wjue7yZ
zrrCD6vDCt1rdmw1AHd5wSkcjJIzXnyZeoX+YYiByP/TA/wHROI4nVsqDWe2c32HntwLvYvM8VDq
MIXBfV8Wr1Ckrtiyldrme50gE21Ju8hpn1Zx3YQSCex+2upB/9r8fxHemfzch8lj/Kt3Iz9Flk/y
enTW5Iju5iPkVPCPYqxuhRxFdHnezqXzzUwGVnfZ00vg9kpr/dRlbsuV7JboJ42GauO/icrCNmom
6mvB52WlWZYCkDGqvLzBQRJsXPk6juqimxMy9L4x+rX/Uqi6lXgkRnnYjiO/G7Nb4Hv16sf21Hik
7MbstuJk1b8uNbjq/oCTEUtZvGUH6kFogFUXB5Vgq9qs2IkR/5XthmTq/EApcCdmgX2PxxTXLEcl
uyjGo2NnB9+y50Pe6SU8vUQN0swLfuiFCYjhRAtL7JsMidJg1b44pQ2GbNC8sKCjzlmje8QTNhPd
xxWuJ0UNo0kD+gbQuOZUt1aaqQbZlubFMlsomX37Bpud1vBeFDYsLRxvYFXTnDnEvbKDW+htzVET
tPA7P3WUGa6Wepn7eZxMo/JG2MFs3Ogy38/rklxsDw01fbXtedNAY1ODtE9eiUrlMjW/PA108Zum
0qJSfnvfT1UTqrWhnZNTjyb3avxLailIzqsDhwTggaa3gH7V5FVY+DPcX3VbOHBq2SSAlHiDmU3f
4BHP1iXeiIKiBNBzCXTMgDYvMqzAQ1nfT0mV4Zc3dH5HMegZNXYYv7oJ5LhXzzwXk+hS0i8siWqL
9079wUYGc19PL7FzKuvnYHk4yzL9ewdQ//jWMBA0znHhKoeu18KqC6rtXTfqI7l8pagg0eYu5KNP
fRaVGnYZjfV6xE2yO3lpZ/JGg1VKA2PllbL5N7/9S7vkEKdpK8nMkkstkhXxRvRsfiRVv3T8JC00
/RCJeGhCtctqddXUFRTfgin/5GyDWGjJDQsxmkad9NR9z0XvoC7uIUSikBmoHuT1/jqGy96X1th/
K6HekLZs61iZA3tatiWAFxlAz7hMVdSLyEzmIfju8sA6AMroG/c5mzksaJJVjfZFB5881yLSAL4D
eQfFqDCnU/OYcikQnVu4WgX9LfDrGiOSRPwzXsU2dIU6evFeJ7kHqRqKk31zupbA6/OuW5aS4EjP
i8tX7FWo5Fh7GAYCyd/H9yYpKnjN6d3S7G1Xo+ObTcZk+HQ3dcrFINWOtRejQVYoOzbDPVnfKoqa
e0zDP/Q5+XEOBPj2fgeoC8GxYzsAeZKBqMBtMGMDBy88Bv86W9TwvfjfLoNC8V7XeFALKTVAqoo/
dHmu3bcIy7UxxCZRk2c6GcKdjoFncn1CDSVZqNLtdlZKDcRx++JsgmqcqMzpEIBVyO4Ikn4+6I7E
ofq6KpCqouIbBbDUGmgJDWxOAyhRp//sVAXLPoKL98AlJtEWG5LkV9LHR409jeg2V1kRNSJf2M//
mzTraup0VMFBnYqVFNEy6iLP+3D0DEl1Ct7JSU5xmIZUXUkZkinyh6v4JGZDh2HVya8MLKVS7ns4
oE5WcZoZTl/1slQxNI6no59eAjqNIGmc6837vgxHl74BAm+25lcJWcM/9zyM3pWont3CSDYN7iWA
/jKejDJn/22kwPw3kE3e9Z3c/Z3MA7K3FL1bJKVfARbnRotjJVmIrz8D/KQJZRVpmtJ/Ok0ZgKuG
DFVKrygiYmY9DBQxvRCYz/yi0bN2+4+x70jH6E8g24fJpnnPisz/LMPUGuJFvlvQqgO0CP7z95Ny
QweGq5cTKdfwgIYCtWbHzB9qqfF3UWTvhwh6PS9AnpFb3nBdd5R8uHcu/0CMgzfq7hBnpYohgqPk
WlozneF9tVpfVCTvCzV53nmXhzWlZ9sGOAkX+5zWKRJjLAcxwShdcme4LA6np0u/xqEVxypgwD6h
8haTMCfm8QsRxIOi1wW12GDlNazuIhZVYWotGH8hdS1AsI3Hw9prVMZeGCQzR7yjrESH4Kc6geNT
Yr80HJ2RtPteoY76sgRXF+JMu2YzmuQkf7W+INPkGw9v4Mrg9JqMLj5LJMkh/8CiL8JBDb/QCDpk
VoGaFyrJqpAwvxJlQiW/woAhkEk204kFh5QSNIMiadZBf6dGiyvGXn1smlFXgg5Azu+Lq9k9SuY4
Te0Hz7OikS9dYZPPv2gwhBlY25Tg/lSLtwRWtgVnqxYoFvH0q+Tq/23iuDnkSHUVg0DhYPdwfTKJ
rDyMclBL47zfTIKihd3Zl1E9cOLAtUHzc7enz/J3B3LeEFP3EWRXYH0DPpdyZCxDQZjJJtMRHnS8
7tvc5yt3xw49wRlVSm7hhRmtZhTxlZYQRuVQB+jOmmGR2DKQNm+9OjxV3wMtPcuPg8oBQrRWchzd
CYK04cYgvCSSNTfkdSlOHOzQ/S63AaNWQmB+PM77IQpRDhPqzM2mmwY36ZfamHl3Azj/LWzqMwpC
VV0bzHWOQluTWq/oMgWC5UxC6VrOypSB0s1e7kQhcHyc5uqXhUHFD/oVLXchsnDeu3ZTYOk6PR4N
YI3trVrTVJjYCnDsuUR3RVMMJ6bVU/Ddiv31HJ1ptTIxtyra5LkcB/du5UWyPyCs1/a9/MRDxs4H
ybmbenkvHQDvkpnHbGNj4A6R8ZVdhW00WlAVrqrT3CXJXiB9MLSsykuTH3WijhZQIRXhLgQOyFru
ZGs7vs+6aFmEfmc3Kz/AKkEiMsvcEuNblIS28gy6RircrXowK7vcWOrA2hht2bdI7/PI7CKHGoQf
kmHHuRlLIyrCCMk/UKISBQfGOXuaRROwzhknOByUO/w/4ClGcocKaEI5QKiwgWJZHykFa7hZZJcR
FrVYhJV48P9kX179FuMTwUXf4Dt/uZL0Ti4b7wLTlsQ7+8usse5cND5wdg79V/HOwWVpd5TjN0pX
CphkorEPC56szxizO6NxaeKMOtyVEgH1oVCmSGjBp6Wr+DRh2srX9lHg5W1OccpzHr99AZBsXtgJ
DqxiDlV79uy8m9OpWxGqQ6cCg1IwVqv83260rD6ZEqXiqesZCulV0zEcnqssxof1sB5G39zjCKRt
bEHDYnSX0wgfWDbYbCE9Ecb5cLzMQXa6UyqPw+biIk4x2dUpIgbv3Epv2kGBBsQe0blYh8gRcIbb
jI/fq8w2iaT5fJWEmjznhw2C3BiEYhLpGecXOuBhoTQyfUulsCxq+Yh/3R+0fUq0ZKWphALwbNvp
rrmdHeby+t/KMqJnRwZtBRDpY9QC/GdAynCtVJTDS3SUob1nGRFnwHchpgNx5pyW3gx9DOUfuH19
A/OWzvM+l+plsDJvCqGxrpfVP5vpXitG+0dk90in+YnTiwbuffEPGGjQ1mDP0fHzw0yoO5YIp79h
Qo+cmufUxgBCRLXJa1nH696mrXfAjc/feXNVk+jSjIMmg/6UV1OJMdwX25QUCBMj16SIPO6BKLZ/
aF5CSdZLqledUIiw2Zwdl3yQ27CIutX3VZVfZK95Uj0RDf3sNJVN760SXjFxNy6hps7SVQbQWS9z
ZKBC2vS1hMq9LYZJt0veLh1YixQRbRra5G6506TVQxLoq2PH7fyOuDXZQMQqQpi+INYwZ+unXYPO
gN1YnsUCMk5FGIFReGqxbuwE508TLsYNlFyPIK0nm/W1eBbmPyqB1pxcX046f1WiXlym9PR9NSen
bFW/owtueW2Yomm75PQ0oyQVl0oYmBmB8Gkgk3vB09aZzqSpvjN1XWDaSeV2qWiTkxfsg5+R6QHC
KkRKubRIbzZf1R1Mx3U/7SK+IRg720uRSNmCG1O1W181COfn9kHOwv41kIJBoS40QtXxuRENnXwc
f6z7FKrQuXuYynZz1KY4aDuCURB2s8rCZ3vyjwUTqMksWXT39yEBVGrWVAbjikjIWL3tbSDg1NSB
BNZJHszf6mokJsMaRON4Pp4/GbUeKbNfrgx76CnjCyxo88WfIZLg+kHK+sdY9+Cdig4bWVZIrat/
4KjwzCj+uwzsr4xSXAmWl+X372LSdLtWUbvWKEL0x661Ec0+LcsPSZaFyjTLYslS++51F6RT/t/D
8gq/5zbNidvFh+Tz2K7kQ92UXSJ8Ml9tfZ787kmBFdrCSebDKd5ucq0VwXDc/nwxhzzAwMhY8lL8
nfRwsCiDEPee/iVV99KTeXTRqJtpI5Y3mGjkIM3tMqmXUEjOo5Hmq9TNpD0UK/Zt/5QV45ZqW9Us
HPP1+0whAX9meOl2ZrG0yomxvYbc2puUMpdHC18zmy2tDDQ+ynmYtwwgVfUzihYc+JYWJ4dhAUAr
ZaeOqK1zXZuvxL/1FRFzmTvNmnA91+52zjrl9jalwgY0SYVlMkFykfi5E6Htlvml/7GpnBUnY7o+
VPDT2qePh654pp/ZWx0JXI2RNULdW/g1VEjG9oADkmMfNMRRqGoJIbo14QSEvQ8WHqAWeGahXe0r
49HJFFjMRI/4XP1/R+pkY8QUmOsn6Pfxh/1ZxYDEf/V4BBUTSpUuEMeSfZM8AI96afJ/GtuG/cZl
NvYTnAkgmrUPKDD2cECuA9HRFbFI5kjBng5YZ4goN8ZooPlDisiJcDe3mhfjA2+DFfsuZOOVd0um
ediLAsWrEctAH5ncn6TMVF+rRTm6Zm37y9M3l6swQ0RAjfkkHuL71zBqi+VjrURkwi4Bn+xcOme7
n56CprxZKTfkoa+uuKbAwnUSdZmuSEqmKbpwpYkFI3yahYDjpxLm/HhzhT/Ur4P2UayqH0zbsybJ
HEv1V+iVP+rHlxjhVPFqA/RgMSazHxrND90Aj/hwxjRA0bHLLNdWQ2A4WPYb/+OrU0qLm7+YjDrH
3+cxgo3JrpDDPHFunNLz16FApvvqbR5+6rZMchVh1IF73xNrCJqhVH+aIrFAvn9eqM6M8Loj8i+i
viMVGRHoQtEC1TPfq519TWv1uTEYjRib81wYIXtCj3//mwoCaVsYHCprzeaSHMiueY9U6fh9/Xnf
7jABIsCZvt2kRZdo9sAgb/xImzvR4deHDC/jmZQI60VoN3zv/DbIpsFn+BFHlGTOWH2oFyvB7lOp
YjeHULc9gEJEI4HJWemJs0BkF/0/ICAk8RcawFva+6GxZQB7Z2TViOiSwJ9HXGtCjYhEGGohHYAu
5QqnYWp+RtNe526HzUj7UR4xMgoamqK9CWya01KzNq0GBy5Uszl8nKzdNWCEvPKyvPQUNmB2egES
vQFS08mgrHN5c+ePe7OJ+iPH9faX5l8Y3NMmqNzrbeoVzDLaQsyOUN2Egy4S7Uo6RF51RZwVjhsy
2OgGGRIiRH4JtwNqwO2JdTTXAuUC4Ku3KbRekWOA5H3p+/7/8cTcUzy3SwdOfRCEMLgG5JG0OjG1
K3ZKITr78Bs+ycTd12p5DU5MqY8eKiEjNlIOVZU82J0nPfHBmPN69BH4ukhthVzMcGUZR6v6N//p
05mfInQC6QzK8WEOztA1glk8WS5caclHuVhnFiwYc5DzcyyYSSrHUemcwL7f3ZaEoJuExD7pSkP2
ggsfTDl9SUy3vfNVyt8ORmsRjEs20SZ2i34J432iTYNt25+NUjzFUQ4Ht5JUjB3qC7pw7ExfjJmB
rmgxiB3IWcn/YaAXqlWxtvuZAEq/psDH+9i65szlwftDdEJyivu6ILueoCt59ue7ZkgdA8ipLVyG
10negCs3NIKrRINKVhOqP3LIxI6zVj6BOvzIe9WWz2zctSqyE6icNx3QLnw713j+oD33L+p1k9OO
q4DEKQp2hlipOIXJI0wvpImJVoPM43ZxDS8QkwMJQ6tWJbdm/F4Cr4ZN88r0JRjUQviyvVKzZypR
funtZQ2xElBIc6edoeBWs62vg0f7T7QurPHVV05WVB3FGlhDU+bi1X7wySDXoLegLpumWoaS1gy3
6xqZ6JlTZKGo0TSIBIej9YV4PukAInL6DFCrMy4WEYYcr+Ace0nCRMTeNkezgcC0Og2uw2UkYQ4U
Bchv7NxtWOIgZuBoI41QBvpULx9RwWy7l/9QijvBM9x5c9LTwiDY50eB3SLLwQImvuSysNSn1oFX
XgZ7AtRXKVBTJEMdbKEnnLSfrY1ezqtaFj1xMhZeL1n7EO+B7iO1HX4CFBbZd7szpYyAd0i090Fp
I62etOnUTVjvCuZu+dzMdIVSACOoUgmGlV7E2zQ4Ekbfh0skr/AsecoAXkx2Ebx5vc0sihYVcO2+
RtkYLRiMyerSYE0eORYuuzsamJlWJWyF373fQOo5nkbnyQkRZ2rX5ZIwMDC13mxaoqbik3t06tH2
NVqp8N574tWytGw6YLLrjDuhFEESZpQSOk0uBAQYMBcX2qHcv93yPiM4zuSxWjn3Ab7ifuh5vlVC
UcOGQYzvWwtVaMn5Zer3qx0kCLA/9Kb3KdKk3JSsxPrOzaJhvdRialOoMgHij+ZjftIb91/05abq
BS5N1MgaBCXtOC3AYsXgUz1A47gWms0kA8XVZI+IDRodwQDftxUiHKAQ7BD4QGlcvUIQjeHtBt51
vFby2MYr6zu3XsfvxwUnPmdP0U3r68K3UkOCCCr+kfIYDYHDnuDIwkPN+NA0JLNL5/tztlqFoKih
5Z98eGTyAEyyEF5T0AmIzQm1Hi3mozdGpUjvu51pRt1u5JJwcAW0BhBkYxguCiLA0JS401V6AM3p
MfnIthRUPL+PKfbxSS9VsfoGLEt4rzvNQ4E9JpwTgdawcGPrb7OotkiUv8VFXWGnbEZQIvDSpTVK
WBCfWM9At2Byh+Mdjh6UkKLFjBZ+Z+k/H/Vorj0Mc2Z+Q4+o7U3Zd2fnkZKClqzBGAEmxGDMIiCA
FHHUorRwSl1xw8uhVngFz3XPTHnnmHG0NB3M1YH8KlxRN8LIzANIlPC/A8sOob0Ek/+opicAnRdB
/t1XUpDUq/SrdD/nUSgPYKKvlXeJ+B3DdcxYVNk2A4Rjt3ZvDcB5L2jMs0N3Pfd1SbpPCDg6+wHX
iXyWfLmjNGibyVVM8jtgRkS2Vedp+/1vb39FDXdtFIzY4+p/A+ZgPmvIZoRw8MZnkBGbptnguHWe
X6BSL6f2ME08ISk7g2nk72OyW4eIeGNhgOPj3BzoS+LszVCJIy8rkCMNNXvbGgZ+A6NRcg/eEpyl
6qHXOMs3L7EU+M5uidO3v/pPAUciu1RBEoU040RkAyAHSYCjKo1IjmvBdoS+lK8WRz+Drh1D+7+a
xGqr9cf4gxD6GWVuG7/O2BGE8U5ofgOf4BQQSEo5+3ySC0fveBoCjfKHZPadH03QfbIDcUB8CGDj
XZONx2y9FXGPz+Bs39mqWAdHMigU2khOI+NhLA7emnSnIqS+Ht69rU0SRQV55WpN1mrILaYK5LAn
nPkMrwR7I3Z9x+8ZYZfGq8RsdWsxGypmgJas06C2muJ26nBOZJRWewM+30s1RQr3Tw9IQzjmTU3U
Cjifp7BFWRMA8sO4Svh9NunWVIX3IvbHWuhtJJ+8JF7RXFggtzTbmgEga5NhF4sst74uEfwodKTk
Xr/aIof3ZCFx/mSmr850EfF34Nnvk0JBdmNLSYw4EahfvTI8jKSQ19npHkFiQgAsfqOEdCT9sPiP
Wsgzd/I0ICTu0PhVqRCBP+L+B0L7Aep6VRbc+/v62ngwaf9WxsrKOZTEF4H1CnF4FnPM31BGtKK/
0EzEmyJorG4M4hkTv7wfKAjsJlMwwZ91eLekYz5Q9KLoRPL047rwNRNsf9/IlYk4uc/SlBCOM3m8
VzjkR5u8hYDZJV+82U4uomNGNa+iOrBPzayr0z817v5H3j4oW3auCbCS+I+qQ8f4TBxVYol2ZfMc
reVbVTPMnCq+pMUnK50PJhy+TIW6mPUiZGAFbr/OQKO8nDXLVaQbnc7sGgp2pEyWtLuCCEdehUEG
9c5bEs+aWV/OxeTIE5rNgdlRnSp7i6hvDmVcKGcsQOhHtrrZt9NukkmEeCUy81iHW/BBoCIKFzPe
r9MeBbenqbWy6XB8L7Ea9vyrHE+w5Zx/femsv5I8hPn0cPvJZb0JTRuV4N7sN7WQ08juzBat2CH0
PMyuFIvy5G1CkFmCfzgx5SdI+VDbnHNH2imfF6mq9DV7E3i0STIVtitruwyJpOZXHZTKUZ/WZ3FY
ITu1tRh//kMk7j5b//+uj71tqAFuRrTESX4mwUTwW+l/Uvwf1T60p1wdEmhKQY9xlJsHOp6xKdH3
K6XkTxWOfq+UlYMSBCxroVfZRtmOJTmesSZ+DrxDaOCYNkv8nT4cVpanfCLXGZZiKntfFbv/H0mT
W9gqFR6c3wZOzZVroWkxUL90fjKjT3cq0/6R+VdRX96P4L4m2MkItn1PpTDQv8g/cAN5zksKX5EE
ul0dcG9ck78a+P9UNeKz8/2tgsXUkxUGluYg2eKks6KsVTIw8R5x6ADyLoEqNLLWHeFJq34lA2B7
3E+XhoUoq3ki1aMX1vm99NJmEuc754o+K6Qci+WH4wF5kTC9dHXbDFl89k50RrKqp4ZF7NqSK1tf
hQ+LSm946mwP5iiwLiZV/ca4uZ0FjYDz8lnXnwKNWw1gXlRgf8OK9lhzTvAv6qmzaZdayYQ7tqVX
SWG6pzfeIpW1o+Q9BD5HQpecsDD43UCYv0CH9fDOAa9tGCFSij6+x8hF8lWc5qr+h3bRyABfY95b
b7mQnlaJ5bz4PPucR2AcLjbNN0TbrstxcF6UBuKR4rC+I1+r9wgT+7w/5PiwP4NENtyC6bwAqsp/
7TrFbPiimv9bJ27EeDn+Ptc2iZvbJisYTaycnFAKg+uYKgTrGhxtd4a1k8PoZf6YiDxaOWtWm+31
f7+tdyOxh33lDBETsJDxbLvoh81hZuOfC5zvynQotvg9G1mP/OTUzkDyCeSsaaCB9PrRxkwfTTsc
VfL2LI/qf20RuvmqxjvXSX3OdN/eHY0YJyysgMd+Ud7uhUktaQQVHsl2kwAaHEMFygRGF2D7oF8f
MOYlGH/KV1UmzfLYz629dY4XFZmTplc1krKKXOrjzwkUC3eSBizH8LmEUk8dWMHDY0lCI6bvUPh8
7RQZue8aSlIWhShnbFYe191KKdyuKn4LJWbX8rVbNxqhOL4XQZUmXlCz2AMymKcuPZLxQdtv7lu3
O5b/kvWNCWtpltGWL5/UkIg5lok4WXTaUDWmKjF7RsHxxU5n9uVr0PAoz1zQR7EFWS+YdsHKnZ3U
bK4y0QAu/f+WqULneznU08HwTz8ACpGr4mVZW9TzGUaAkY633JCNHy/8xtz0qcxLPSyK8i/b9fz0
808mHD0vAyCs0Ss/Xwi17BX/N5jbsFwdshg3t7FPOcFZAJSfSxmbFdixabP4PP9+fqPBfcz7GoSL
ypNiae5BQGExgZP5VpYRa49hY/c2iU0jEVN1pYGgQAbBxtDiO7GxcvyouCsg6WaX1a5zKmIVpOin
m54FjotoL/XH+U5KeXejIxMvopNGx6Z3wYZi7g+DoU+IlTmNMTea2VnPYlu3qjb08WhK/ZVuJUPD
hWyniEzIr5hh8vWQQVVPrennrvrdMl8OTnPPNw1rqZV1g4JdIsEN7ON7BQrYnhYY5CId9gBpnkhs
gIUsrI2qXRG4irnT5mcMJUFTMNaMBmXH+bzBOvd4vEsDmO+uVGzxKqf+i0OOoy3/7HyEUCZNriXs
DPOv4EP4e3lkixbAIqfiT8M/R6O7b1ORVQRZjLK1qbHoiGQ1HM7W9oJvVM2YLZEnfCBqB6OuqA2j
SK68lxlSFzIyE3YBR02HJ7eX+0RNV4XpyPtmXd8VwmcYY0S+aDIwQE2oNBfk7k8wP8wvBHsWVhnU
V6bsp9nGIoX7YexAFW/CTj/hCVzRlsinSRdri7w3mjKxECfFD9sArvmDHVDnrbuiQ5S5R8a1bbdN
FGsDbo4JK3Z4ORFLap+CkTcgfr1IvnFOOgL+CZNKQFloD65KBP+WLcq+FG6QxdeoqbMNWYU3lvQB
d8FL+7Rrxt87huVG7GecF2X7RQZRP3AU22YFb2BDE+Qw8JHLBTE1SHc5UU0jd8+5tAkSp1Jm2lat
bxlA5zBJm6i7VvQrkvTrZQa43SRxqe/vcN/oPl4S5agS4mAGdTQWKHEMskHxg01QUOuhR3udd0Kt
7uigTYdzLxVjP1G/JFDBeGKrqb/dd8/8ps1oN3GtfKey2aB4EBsTQ7s3lG80oBzxNAR366qAizhT
mwgrIe/MHPKOfTJyK+jWkioXo5A3A0KGC8Ao5T6vSmkxB9J53yv7GS/tCGPZE9dnClxAKIzR+AjC
yOHes7y1m5Eb+q2ndGXdsvLUFNJzJMIJFYvPv4x0VI5Fz6kV/epzZaBJNWov4CHDpdgq2OR+/J2o
njLGF+TXO8zgCwsAap6jlbcj5inkQ/yhTluisouBnemtco9/z1SSOnCm1ndAaNClN2zs4u7NTZ31
b3jc0DdVbmyaFSgZ3J33uZKRABhfijbDRSxkJR28iEEpSTM5GDH8jfB2LFl3oORdMaWMFgWN1ATm
AGrCNTtZF0jUSFL3txmNr/0Tb6DXAokf0vBPXdx/lqeE9RM8sfgudrhyBF1SYlC6mfGhg43yEmuN
lhjZgKq+Q3M/NMispKrBzcmbrSVSOgqxFTC3JjERelnpOyM8xEk8HylognKpo3cha1ckiaQtAYSX
5msRtmbceh+Zw9CXSMek0L/8hLwM+c7b7bcSOfsVopxMIE3wLdMHgd4lvpYoa4U7WGVI634+A0X6
jDPyIXa27dTO/p7UvJOos0a3er59MzeNRZziXbHZ111eyIGLg44CXD2DwYkttd5tqToR+k9NRng9
fQe29FtYwL0u20haW0ssYEfTGGrZ6gZdbJYm5aj9O9YOh4lP/lUTOWkj6+qrwwaZwVDHP+oWnTBV
NRDOszMDG0WsvT89HxxEZq49BCdutYQc+3k+hRPV17yeelft5GdB5IDbqy/2xL806khnKrtMY5wf
YCUpfutN+rgwKkB2CaeLpEJUucvTluQw2m13INHVSYVZRLr+FzvsiO+Fa8owFUoYuM267ky/Vv6X
bEteJ0hzOFm5VvlWTFTBCc09tuBmPbDRuheWt6H1+A3ww5BANDDp1BHsMMkR/kszs+1AFiJvDsgR
uclPClF90gZCl3CIa3I/jSo7TarP5v4615KpatnlPmDSr8MqdvUi88B5Yrso6OZDQU+9qWtseFUk
kiWO6kCuYea14eKG/uAvtzMT4aWqv9OBzD5P7Jp8SpPSJjy/vV62YQuPyPTgLYV/lM+KozU0o8Pz
Biqcu/yEG+mHHhKoKV71gGTV2w50LDJLrxj1OBsJRqZwX9tLCNLDJ76UHKPELnIVCnlZvHodPX3D
7WSo42T0n9QT/vQJ+py1rQaExJDfxxN9xTI0EvAzZ8eaiY9qDlHR5AxdPu9aTkKeEFvh2RuzuYPt
uADTaNFO8vk1m8SomqUfOzTy8m0VAPkQF9nzKFMfL8612NEPqQv8OexduNNC1BzBrInhsbBF82Lt
NLIRiaX74E8eHwVDDqXpPdr9KjMRDdI5Huekz89FWWjmKKdBrP9wtCHrMHsabhx9TYTTr0Lxo049
IE6woYS6OG89lj1Kz/YRTwcUiPk8zyrB549aUbN0uRQkUndZwD37sdAmXwy3JKX3Ur4NHqCC+R/P
+TapqaEwQN3lHrzYhWu0T1zbB2sJ9OXHlif2Ob/hKHvZqAcU0xMVzDypj14hngWZEiXrHfzycBpH
vZ27f62s4ABf6WxXa6ymQBVFH6Dfz1cVgsdUaYPsJeKlvA7duixMkoVtFNcw4oVoqQZYfXNvrqIY
rjkYUKFtzg5WSbjGRjZZ7686fHpmkK5JkcZv1skBsgxqtRpfW9mq2Wp2Cvgg/AXyBdzOunwMzIPO
LQIjgfOIG4n3CzHVY4xs5vkSpl6QzNEKE5eXs5Hr/KD+F09i9Fym5EYk96qyj+TloNsqnL+8+PJV
LcqqZr+7Y4SiVVqtBNTjeUIC5wQnh93mru7iAR2hNEBxh7fh2r/Iij1s+7/1Y56inAZNhn/bkkHS
ScMFJoAIfv3BYrYj222T8AAuHqL+zglap2H2lFWS+m0upr/eOYtBnsHnn4msIIF+DweOZS1t51vP
yVD5opieQo/jLYgZPbcZU+4eUSTO3068GPf3TAERZjDrRYI2H6LgVvHU0jWd7P3AUEFM2W6OZdRz
4fC774jcAKC+iieTyXDyA7d9YvRKpifchUIvBnn7x3WLtOqHAj8RsjOf5/gTLD3wPKmKpHZrDHT4
3cBzaydISafyCFdrPGhGqAEfvOGxZUhfYlh/Z97GId1PrwXY0qKsXWS6DQuhLKKXuoxdS0uMzeaM
0TjQbfOSmP377Jw5ajn3deoUZsg+gxJ3/ymXGwgrPre56tIu0dzmSbrx8juvY0iG4sMBZs7KunkA
AoEEHTGJNQZhTj09EBMgIv+f46cvIpD+azmeONIhZTlhkq33j6UiesreWlHhsNL7qF4nL0C1vr/F
7PJ5Spr81Fpub2KcUX8z8y26i59n7cgTPwDlIk0j8jXx82BQ/onsUWZd2eCNn1MBIcA9L0BWy3rX
hYakFXmx3JtKcLSm/sZ8owemTs2Hd51a2qe6E15roebBvJhf3ss2i1pJZgCN1cleFJhQfZTkDc/V
vrKaotRGbZgagO9Urckwg81FtDXTd8H+sNE85EuqrFHrRQivImoG+b9jQqspZ90hN15sGUY+rzP0
ufqlCUhNwUu2bO+hdC/FB2K54JR8kAvUY2xSdTsVtu8iOXRO18Wz75h/KDojHFotjrhTqKJD2+o8
XMXFddJ6GQUbouBI7nAPFjLIOCYV5gOV1QriK3T+OzCUIY66oSwU/FxpEh8IZNKmSrhP02X4mnof
icTl13ycTxruTnetPcrqPLRP8QMED3smuxl5fgCwwXDOkI9B+0axwmDJCudPdX+Sdafm/ugGmQbd
m6i0aHyz7dOIAaHz/YZHIlsrL8o7ZuBFs/MNIlkVokuRCZ2ZGlXVyA8owZlEd8T/d4S8TEk3eosD
nS+O7sS2lh3Hwuso94N+qnJK8seAle7CaivAQLgd8WiKTYzbfoEg5pyY/oELG/BLf2JnPVoNuBiE
al4YKvLI31YWpB2tokI14uQskWkY3HeNMSa8MO4ej74PqdgfudU6qVY1ZeU0vQSd4Zbp+KJatyXQ
tn1NcLrMzjadXU6/BSbUz0nzdhZ9B6/fn4EL76GvMbCzhAaHJ6fj0E++8qDyTTaJo6QwW9ZD5oKC
+lU6vjN3dnGmFUgFEvKaTj/a3pxtCNJe+NS6NB+P/CNtTqGykq8ThqbtRbLivOQvZK6SH0poRkGl
pXg90cQtSkL+W/HaZknGo43v7+bhrtTVm1iHpkTC0o7/xKMCPrQkmadXtsyvvpuyOk7TzGNZhwfu
/O2RfXB1NTQy+FEvZObXg0NCEcF8q0a27IAcI5rdJ+i1RuX3mNJekvfCvZV6xtuXX5nKzZiD0DGK
pqqlDfCZMF7j0qDgXHttAzsSJlyDs8sJKOD9TDGX0T1JCVs4gxecBznhrBFxkujAFHNIf0cLJpWc
Du9tugYRBjVfN08KxGNU2wiLhPHA63Ol18dyWOztmnlmVkFmWrsJd1QX40dSjPYks/qLHE4s2ulX
ZGvP213O3ljoj9ypcmk2VSm4Ztvqlz1RSjcXG02q1SQZtHkO345dyvO2dkF1rNPVSvV1gjVcEBOW
jl+3ARBTDnM3HI7fgckFSyfyr4v0FirWVannxcyOUE9XcIxltDJupRyDzePlMhkfdf5wWZkOJYwr
tgDvaaFBFaasbgvLy4vdn8no8scB5C2aGyEAOF1/0GzEyVy5afq6G2sWEVBLeHXlnYH9ODeS+DmI
mI3WkPCH7q/WHEI32BbfjuDzY0kOhYNsRhN0bLV1DvejdLLkzQadJJ/THspF3Cp2ncS5vjQopcNV
D86vm5rvcXGjZE26Nt7C3HaStLg8xXGwlh4jqf9i4TCQAMlmOqQgzxfQpGBLo29RvQfRlIr225o5
irSQrjxYpC+ammFD1o6CNYSpTCM2Xe134AEbtYSY+0pGHwoXvqbb2Ir0/33qhjf25uftAx2PPybZ
CfKsJND80dfaqcCVMgz1/sM5nSW5W046b0PjNAxYDwfEGkiB5I9BmDfr4eN48nj9YbFHKDSlUxJd
tZY5XM0WYuAoBpoeL7LlVBK9sP3dO9qbezAjubrEapoceK24pD63o7l8Kd+aIeGnJdjwk7k/OqRO
/161Y6s/BEzbjWt8XUaHdV331FiWFqivcibrRgai4uYPBqF575F1pxcqSyNYhXXQXsD2QLx1LPC6
AEI72jIO+Dyn7OCgvmlXDkE7FK4nv0UqoV72txsXdmkjdC19qOgOJHW+hqaVnxDaKmPmc6zo23qi
TJ3ewLzPBO1h9NqzGOAzvwIPg2l1oM1c67Flg0bffLTOZ5uwhkponnKqDs8wuheN9wufBIb2q5Rf
cK9XCuxsK2779KpYdAik7ca7eGcABooSLSQm1Bzy7xLOoUWKBbbS1Rn11+LeSvPs5Iww52CHjV+S
wS5+Vk8Oq7Mh4WfYtbj9JVTwJDNCi/ufq7ZnKQFKw9iNc7ZrxRHOtf1Fjx0If2J9up5j/o+ab9oC
DNcDyOOzOHTtPRqdCoY0TvMIV6M9YxkcGuFKL28p7KrEiXp5aYL/1QCCkhdWzfo7aKoztdT0F6Tz
Ib2oJyzrA8rGBhd3SkeumOcoVVwBMB9eh7lhduP0P9qkcMANFPzPWPS7ORjdzDdmvNZKsYoJVsl+
YIb1Vm5tAc2tq+PNalhibU28HhzntQOhJtY7w1E7wN3G4L2gHJbw1OEwkLKjeBjEr5CUgzzNrRdJ
E1FUDVRIigi1t726bXMReHoHXQ1h29ZlQK1x5OZRLlqaHYL8d0HHgy4Un3aCR/JJCZToDqRq+1m6
1kBSwMo6WqxlFwTUuEXkysw46Qlut8IeWCX10YiIGlbjvlOwNViVBfEEj15cDZONuMct0oUrmxGc
91xEfNA4yPobMXCITV0G7pMt/bTRyFaaD1dVl7KQueMqmtjeZlN8NVFq/zkW2y9vPSUeYgAtVDr0
VM8HpBRYScoDo7WeCi7Pc/50DZSu5Do/TlvaSoSLYWUe/J4R+Uj6/ykIE10M+S5H+U0itTEqKGX7
91AHrQcQqOJeHCGVVLgw3WtRPUeAQbWpk/0ouWKm9Nhob7unD1ZJwhZJ0pF+NVuRVO1vm6P9uhrx
TL5nEKM79U4eZ2KhF1F3eEbADHChCfnZ3OLzyQ2hyC3V+BAVQo2Qq5PW56Na5kNPu8w6AuhOWgnL
hT+mBlkEfgR1aGYWW0d0KzFO6ckTLO9Vh1q1Tm6+05x6vYdaFAFHcqZG064OjiG4l053kC6j4Ngn
Ens0ZZNlR4cSe2aixV9irQi7yXJqmbt/E2ck7qTwXh55D+elwXV/J0zb49RuPAD381nti1HBnMc3
OZyolfzAIap23f4oqMPHkTLqPu/M/X84T2sQbonN7xGxI9aoDw8+5dOljX5vPUrB1Lm0OqSHhhOw
kulyBWkQhDsbH7LoCZw4pVADhjXuJzsOH1+8mn8NHLtd6Q+GtrgRVLcbvd5lY1bFMu6Et2LcIA3V
6PTKa3j/kWHvT9NpiaE6r8gt2XnebhhEg3pYVyH3d26ZVs8bbt6n2PcybrSZXv/uo2UM3C/oWksl
35+E/ZEXrC2uHXs2xgEQQ7IWhl8TEEZKBBxHIo4OrWWrAqnuu31W/QCwNm8wNlDwyGtZ9asHa1pv
FawhEQ9gQSzQQRCVDn/FKQGnrYBosAUd06JGGnafUalHgafA7Kb49c9DkGZ4AHzop/0GUQT+6r+o
iHKZm5bUlefnwr6MGgxPtwYlgNpJfnjLWqtMa4aT968pR84U8nLajfD+HVrpq3qYUUYUQfMPCJ8U
K6xyz4y2+Ewr3y/uJEZM7zjo6YbaKbQegipLAz2veugOQrYsYayUCGniklVWn5rO6HxEqtALO0OC
6ZRkbq9XkjeOFdv6xvXL4bzUNp3h+h/4BQLbpbZFvy1/wiPPnDn/4zUZLUvPQ9obh+hvBeCKwnWH
0xPVK5FODWbRNDBmmg6MmcTBRqg/wPniVn/oY62ge7lOLBqJ1S/JLfzLC2T1A40NRl3kGWnP5UdZ
QW3XL4DoYxWeNl0zzhlgh4o41AUHJcXP+T4g8WKLYSKbvJTMHzeXiYyGggXfJYhL+yoZZQMRuHGm
af4L42s2z7JNV3Z+8TbXqT6puWp8cjGs+Hu6tT0xMErguCgxfha874AyKmrlntz4g0L3zqjqBVAg
s8Izi9ymj4D0KXVlvRsZIvUmxxKO8tUOG+Limy2WCiAQFgRavPzU7OwMI4zu08xMZ0S4mTXj08IU
LYK07g2L3EpLrwdWX74JAI0q9lnUL/JFLZueetcSU4P3LSKwNGuDQhMTT0d16RUx0acHgOByAPLQ
aN8Ackc7EkJUP3jWRlRgyFJERwJO/o4n8o32/vtrhnCtum/jxFNXS4Vyv9T2oEKttWDAlZSreRUk
bnKR/9EJfr60ouVlQA6ADtp60LjVCAeJ9TZH6FRFuJhno8pE9pqk4sl3m+MHQ3jZPJ0i+1J+BRT+
Z/XjgpHacBMVkeud1FoZcrMpSKAMf9FdKzllweYGC4R+NVwZoywNw3RUbiEskZFs143vjPFccA0O
BHYBnA/D9uJBOQPl/ZMjB8VikCrjCc+WWO6onhnVBIevY3/ur2fIRffQsR6D7lTGYyfEOo/sOEAf
fw60S+1v9NlR1KJuREdQMGvALSXyNgdVcnIRktMFCPp4Fs3C57jUfc8cES/75sWq/70EpBe1v/9k
G4pI4mak5HMN2LXKNS2gZGaotuJiaVZswK/9nZo4kdLPoF5AKYTGFnc5fZhmXTrYnffNRGDz4aRX
xt5UWEyg/NJnYdt/hnjInV3hLDpUgKdTdL7EOx/fRICXJeOND4WZNXFAXd3BOjFsJmQcMpolmSbG
60zgckR9+Yn+l0NlF58xFxFRrIZqRWXmMxA31MPqkE2LXL4x2KocGeFsKKxgy4807CL9R3eytrQQ
PBoMcxjElvhyp5WCw9AhVx9OoDWnTcVsbtgD3VR5xKuQeHmMadUVB9tmjNc7YigewUfAvJMdIGrf
IxDyyNQPu6JEbFoDwrX5ArRWzfKehbtn9RuvvrGu7rv69lwWozb7i++wroBHZddXVnSAmoT9wr1E
jjCCr0L5y3WNBfgO66mPsBhoZyuyzPjx62YbDA2Z8WGhjHVGMqXb+B9Eepyb+FL0qqKI56l4GE23
nLiFJoC7nXC+0WnlQXVCFKpUwcr+6g8Ccrtp/G65EB8M2pNpO/04qrXmiwI4Kqqn0RZv5WdYsmko
P70hFG43ipbgJ/ACnuvpqrHJ1Sevy4oNk8nDYPGzgtD35RD5evkLSp92TBxBrXmaV4v4BtuuBw8w
jfwxFGsMLk12N2ssFefVVUKEq5Qi9UEJqofYnTpzn8JctIP/3O8nbMq0HwTn3RPFVgQvC5nXJs6s
FwI9eWWCeV5E53cdtil95NNITEuUiOsJ+9c3s4qK/0BtgTyPKs96ZvwXlyU1ecpyVz2tFsX1eomS
RU8ObW8BZqNL9w4T2ADZaroTz7ajXyta1a5+nd0IhAH3+c2n0z4JYEc8rdVlgD8eZ1h3xtq7Lh1q
LHTuUTKU6asdWsSHUNLy/WcOWRXCPEgos1QopI2TTBaXukG/2B1sOmkmpSVJPIv9g+h9bgS8V/F/
5ATvivyhwtbuWFSwFPrmcdaHAP6gcAYTlV62C6yq954auSzykDGlWZ4z833VH0kHrmBl90NvujZY
3Kacg8rijB6tniVS8cjY2MXkXYj/LIVoc9sF4VvfSfTcjyIOPoB7/zde0xYRptC4O1k5uze4cR3V
NPaYiXn2m9n72ekOrIOwne/MiV+HLNWqzSLI9TrGJZMDnm1UrxU9yW5/qFlLUkx0Q7yjFC06kb3h
HLCvF/WDuxUjSu78G9f4Rwo12y8pMlBqgcsM1rPGwsdVqB3GVeLfCWsWDDced+JRG3bH2cZtsMsC
HYI0nka6LPN71Eba/fXkKP5AHvBW2jgLq8PQfuvvhAn49ONz9Ns1kIXLu+aKE2QykaLM+zGGRwoK
LSsS0PhKg3OsAHyWa67m1lPFbk0uHRCHZkUCSjbAqDLHvkkC1CHkxik1rMdkPbQbPon37tMh4Shb
+MieS1HtjJcE2AT3tM/AF3FC8/NTuHWks/EwRo8suc20e7mvRhWHhXWJHQm3ELRb5ZClJqguy9PI
WC1uZ7znimJfTArtMJF6eD2OFgWIqurmNIelP0VFLmXo2WQRXhej+DT+4aB8GcOjhWOV1rlVez9o
ReoR4zdWOp88xm+vjEa5ugNXx959DpOW78/x9Dr3URmGQm/uDt9ib5dA+dOg3KhnQHFJIsXqNoWS
bdUZ053coVUewQuh4V2zVo4pMd2ST18cudNAwE4ZiKhg8PKkuhwO/tKckrS/PNAjtkdnJTzzl4CB
uoPe8I9Ou9yKiXLidvTcBON+Pp69JDXQ5Bh9N9h210SWUNuOGFZ5JWzgCTa48xnzWEdjXuIaRU34
oDxXdtsELq0vRvwYtmOxSDgDHMwp1qlm8UEobqQtgDeUyYZPrkHGo8C+zsl6od2onldqp+yBDob8
Haj0fDV0vbKNoQN1BdFBmOSeLTmWjRGVcik0lShG3277Wn4n6cFwmxH3K3ClG44gwyVYhrCQ55dX
Qxp7qGsBWIAi1zIJ/enyBF86CNrK/Yl39jQAADyJ53UGFAEvPMfVzI22yrQHwnE/3GfGh/tHDeDI
FKQqzDEWy5YFtxdjI500VOkLAiipZGAAoF+atuAtZrgAQCr28h+WtoNhKNcfe2K9FlNi027GMEhK
3aOefxaprWFHGl6VUD1hKTJDr6/1KeNZptelBphPTufFU2IJHanaOA9tGlycuPH7P8DrZlFHasxn
tazQWnG9wB5w1ZML5xXuhTTyi7Jl42ks39WkNgDvtufGaXOq503FFvhlM4AxiDhQi5HwCIdfG2Qc
J4H5bGeaYwTebWbG5FDtwZa+vfuVWQ8g+t/qKpLyZxrZyLna7eU/5XsizL4Ga4kig475EQv/3exs
0MXUvXrDnCJ4xRZ4TG/31bJFg2SWDW3dtYJbf6dYJ4tNnv6xK/9moNyEGht6Z/hT0AwbWGIqdDey
XA14mAU9l4pQziENdfWE0IWq2tkaqLJTcwmxayQ+nH9kcTiXwbyTC0+Qx7NEG8/Z0JKyoAAGB7Zm
fKlUR3dP8HaXGMOefMjTEHq4DhM2YLfzKNOAGiM4SOYZMXBTCywn2T4wrZZlB8fg/VV3smiOJSW0
GL+OZidvyfoF55+hfezvr38lD3O3g4p+j6xpNf9/R+ORHmaFHrhwrh2J7+MhfeFfB8HG39tedAOT
3gN4CBzno3+rbZ3yR6GeXBDYEf6qtqwjJTgpdHdbWmYy0lx7EqmrE5lskL7NHy+POP9xWKlY5yQ+
0zXpBVYhJmoEF03M7QTdXV9g50iOEY83jhThogI7WyOeXD1FjwArJ4OzfZyPnkti3oTbNvkJ8Ur0
yzCDcvetYqkGCyr4ULqmvQPMLx/5F9zAC/WjYpnFZuwd/qfIstJVIwMG7GRvVpJPy40RwQyAN0Hw
AsVp4l3WvBbhaTzCeVTNYxB1r/iPRZIgp1p5tljrLQ9E0z2kBH2K834heC4CJyQ2zkHT5Tf7edre
5doOPjqXXyoa93hL1g0cEni/uFinKCNw4oA2/yvZGMKl38vd1ldOaGptT1xLS7m//r+9CKV+sTtV
0FfXeSUo8wdAJjRySSCItVSfc4P4r8CP01qINUPkci2XUMhzvUSFeX6QGw6gzL/zuQ8Oz99yUluD
BtM5rYI4RfwCJFYFIRv7ye1tFxD/uqmo4QCg5ZDqF1aLbhgKI6MxbbAH3SDm/WExWp3a4lUI4s9l
Q7wUUo24xOrfBNjBgWho3HVWNLiYFrlOFomQporB6Vb44w+/5GZjeVoXJIqZylufu3xuvB2nsq7u
Y4/2gE4Qzsd0BktuQQRQMfjCKJPjhlbArJzgE4lnJAn7heqLgXasoZS9U94w5BK1QybD2MtsaU7s
y+OSbWnLXiAGaADZBZPdp5VT0bsFYxPNe0gpZZ/4DeUgT2/lwUfh64StQ4VcJ2eFxhTRaPRngWYg
9JPjCqBZ48iFTQYOjnjmLFSxqWdVLvCCa7BDjcDAl78E8RWWf6fGBskIW6KlaCokHpP8AWo0BiWR
diAYVLE8OFLnsIYA3v8JjYJGUrijY3HcT4P/d/zjXKri4mKenJOQQVB7zwUpBrT5yEZI54JKN+fG
4c4SHwXUWDvH9UTvJN/DvgCAo2erXuzx7ItdejF+uFnjkvo8hjsHMvHBogdC4Augg/20yVLk0djE
WhxoZiM0JXjj5+yNFgPwkTHIgpL5Bfamdtb8HaPVRMyx7AvR/sCH6QVwewSnAI+9xK3sfUorNx1V
4a6bkgKhfKtKJ/3BstChQPMO4rdRwGwHTywQQfzCN++JQiEgXIRBOaygxSQ4zS/4XAjo12/CXty7
67v9FFGviE1lnpR8uC4dPtWzw6g0zKGcNFrnFMZU/r3RRrugZzoTbGkjSX5049Y1oFKBRhndSgAk
64T3v96l1yi2uVBl2dAJmfxoh24SSFvG82NMysIJjG8zCKQ9N2gW+zXerM3WG26p6chEfPYuGb67
M7Ug1FfA6lWPuwiOla5DP+1IpGjYIopzdWJqGzQplrDXNFoceNeDBtpSUpOlcyEXsZRBk6VLZi1f
68THbYOE3CiINVvUL6YBgewEY1dZ8qKq4wn85rSW67OFgfPLjpkTwmV4t9aVy9Pe3vwJkFLoxQML
4oGfSFIbMKCzNsG9oUlZxXuQvZvcUB1AH1Q6uyzVVb6T7R1pxqYhbAKAo7z4Q5ieMwKfhQ1t6Gg9
DjXdy8YO3J3Cf+Z0dcn8fp0TPXSfSUlNeDE5fKx/2s67LkTAkCYsAQohBzXtqUqIRz4f9Bs2iRJK
erZQHPPzZznMKHrgWJS+TmcE05ERfjP4wKxE2DYYZlP1KyGM09Gzl9ajnXcjWP/JkhN8H4LCCwFZ
zCGpbYWQjAoNDk0yINlxbAQVeBLY8TgVZ9a3Gah/T9u0Q6n60UWW+oTY7aaBrx6zXs0EfW2DkavW
cFd4cdSd+uI7eWpTLiSsHbmk78IwUwQNJNLjNYAiyH0WtfH0GZ4+hSeh/l5bINfgfEzqiLz7KI9O
0pndI2V9AxYKX/hQ30NAR8yVGMuEaMw1XevrLAuBZJTkdAviZruqkgvMfYWCsZXcR8bb4VZRhSc7
zM+v2Uh2KS/SIFgXfFjJnvgeTq/ERBJvIe2EvWbqgmo293aO7DHRZ1Gk29ieHdMBVnQGrOgRizUA
4Pby2waZEXmRLSSVfzzw5MPcxmoV4FJwc9TYAZg2AEULJ3rrNCZGd3Y1VtgKF58zLk3vswnbBIQp
N95pZ3ucrvQJoppo9EPFSXeP3Kcys52SJnkFhEZsm57PMeCagunvv02VaS6YqOOnN0MCPfKupxG8
ag8xcDLSj3O9R6rj+vwjIaOkdvUg4CG+6fRy81uzawig/8vS3q3k3DF+L+OIk1kDeS/RtlgHxxxx
jftGPj+og9GzJkN9hfizWjWHeuE7aqkaOKtexDqcIghJQea+zUuB4xjShL43ZyQo1gRxApcxOYpI
ip0E+mALEpdIRhfGkj35myHcsbTib0uG05ANScPDFK/5MV0R3aojLLN/2D0HP535ZL5Tu/y0Gdrj
VdqnVnek5oNSEczlRTJOt5IvPsmu/Wb6sPAFK9rp5xdgpxhUQudeNgCzzN1LKZO2MrPN201+jH37
9nojQG8lkZ0b1Bj07nihySzSxOxlXHRdqzHw664+jIdF5I+TNd2CVQCEy5yC91kGkJLEptEwhpsE
Qjo1fNUxfegGfU2CseeGRNHT84UmWDPiezyMJrYKURu41cNdOnp0XR0e5GOwJz8l8/UGivoaKWxa
tQaUPW+uumLHA8cHfqJIEzpQfB3V5HNXcOmyiffol3JXO5qdHnQcOICikYfWMF3TpuZcBSzGGrgY
COfRCw2Jla4n7QgA+N6jlQ5gSQ8JQ2n+12OVa3jIx+0ylPadMYo7pRZw1/IW7zBMoYofZXaexXcn
MnrKYfaUrPllQYPPvuvW89KJrjFIHexAQ1ptYDNghymaHo3YmIKGqp/NoI2HI6VL6H7IARwfshKX
KnZ7BIyFpPIB3pTwkVY9wKsvXBUUtTq8YiXjzgbWDB/zn1OwHR5H2OaMM9wLq4Hq0o8Qp6ShdLe0
BM0lRuNyWEn5Ytu7rn9LhaqJ8P/O3W44HRTLs8GHEDtkt+CNRoTgbP+B6pM5FNFcAvvYTasJ0Xmd
EpmD5/BMc474Rw8y1ctF/KWRvDT4inclwAHgo/Ee2ZzpEWYwkOgRuausA+L0lNflIKAR3/zBtsoZ
VNHikWpZ40eS5UELoKfq2IY1Qa8yhReNJPioWhN1bNyxZ9f4S1cb65FGpcZ9rtxlXWMVO56c4uis
4nEdUl6I+xiqNscdU9VEAcQioGFOAVkQB3bOnUmLQP7k0diVoD34kUkCZEGs9IpSlZ4FZmRruexx
aqw8GOv4bPD5mDWX4OXZZrdI+EdnZTQkeo+s7AvSrl8T+oIlW56o5YcHt3SLtRhghWcwkjMLaEcV
DoOrfN6Fwtmr5Enosp6hdCV77sPngiBCzds+duOTExJYX8v3BflJSr4hA4khgrQOt4cTuhh0efWs
1vdaflSa2AiTtv3wNmhA/vlRA9o44aaLvDi8cDuV7a0hBEELo/0xBTlSJbiLOXkx6a0GtCRY8Dfz
Qx94mGtnPuk3Z4IdAzMIcVYny5J8yUeLHlAHZPnUiuu/g9a4+epte56bZFUFOMzdN/rxXtAj13O9
zOx0/RcDtU51LH9BtcLMebFBC//Y80bVvf9jsnk1h+wZPqd13ymmrvuVfFoCEcKXSIA2Mou/xjIN
fwi4jxUI8RV7Uff3nbcp08glpwPeCOKBHDcbAzzjf923dyVdNEJrKufQWxFuhEy6qLcXNSA+sZta
iWond7UhUQy9kIFsZiWNn8iHmXKyvF5B0EukasHJW8e59jncwe13SF+7mqHvJkTApKRy8Hv5LUfi
5a1hU4/iy2+6rxUluN4tdJTWfQpQKa2YjUaxyclEiOuWpantp/scfS3gl3tlv4jhFsRd1bsNQOIh
+nGCAZo6D9MrzsNuKtbTwD3krKVvv+VNb7u/8ME1SoyHJs1890rk+2X5D9iRe+gac3CBM8lILsE0
ZrsGBbl9jMMUD3eeY30Mg3QdgIKHw1WGAgt2LyR7x2EODbywjuGayFSPtORMRSq1iK+htYFvSwHg
0FxXN8YPr+IF8TfzZv3ZVkJUppidqIR4N4Ke3UBmWdVJ24yB5wcXLyNhWpMWuWojZyxUG9M2yIt4
JTHNmxokrPFLSD0rt4eM0ahlD/8aUhmYAJryPw4pSr00fw8hL5r6x+hJ3dnZ64C0BQBhP6oQQyX8
2Xpv448tsO7LV+85cclh7vPXiDx5pI0wzGUYzmsiv9UaoWsbjMl77tTXcWovXVoZQsCPXv82zhwu
r9UjufjgHoqXMMXLkxOhzdnlVvWAYpjBi6hqUXfl6M20r5K4FRtc0Z9Gr1nmFLvIq12gzYX9l9yb
uVACnWt2MAeP7L/kX8yDv3t7fru1vIV6Nn0bEDIRu6arUfvjlsZSO6xNRVrg2Kv6i+R073rIc32M
EOH4dG1FZSdo++In93GIeyiHLcE44fMrEVDQULCABz1U3RlJtV3x/1xJxnD40adL/POI0INLd6LQ
by5EuwoCjgc9J3DEc+uIfZpEEJeEp2u1idQXikGzDmTr9M5ti5MluKZr/sHT32HekCGbmfRbYZGr
TVajrzbB5IUxM+rRfscmz3rk/yH/KOSGKYsZAs3MCBXuQQm6wVg3nqV9I7HQezhxZzzTJEUFq2Fm
cva0gL8KIyMeSbc2269hUtHFoj0O7USR/UK4n2Re43r1TZMvDb/ZFmrCVrLd4nZmstwSpRYSr9bh
dJWgJlfYejp4EZklhyJBqchft4ToQliB3sGe5o/E2k9TPNal84cwShd1mESpkS0dSgmfkutJENaC
DREfRSHZoxV1raXZffXl6e/ZJAshzSfkV/1vdYVbXM7H4ay8L/ggexjiwLuTNeaWk3/a8dYHDzzh
OXEgEwWmoyuCt9bUxuJ8YZVy193+Qnw6TDdYWIkwQ3//xtSAaoLsdwCI/x7pQurQyaDpBH9s1wqX
GwSJDS8ORv1gVRJlDBWF+ac31mJ3HG4AWUFU5o3A4SwapsJlIoWX/SSudtxfVLuC4rAqLuX7x2n+
rbqbRdXTwNLyVVyY2h9st7Na6Vdyf+2qT2+IwVeFncHHiKFd+UrPPhetb8obpxh6qH8xXFLVdLqI
/ue2JE/+/tvO8FDs/6SPBodhR34GdG+Qaz2psSSw/5G7vG8fh1PgDZ1bbSh9YZlquAY70g+1Lxrj
lpY56bNtab/hBqm7kzu57q/FvD07NtGzwNeSW1V3vdk4wIsK2bPtczQPAwnPxsxl3S2ZX4fRie7V
6VLlY8HHDCAa0IbHgmMVbd6P1QCs5nbhNv/CdI/71p9HknH7Npa0H+mjbo1Z9mwqotxr14NUu1oe
nTFcvwGOw3bLKcFT1eosr40zxQdVZIaUgQsRzvj7EDxBrq79ary1BlnCTzBJICCZe5ImdhrChVHL
Q6oQkCUeUXpjso+48K0J18ZTU6PlYIIDV2SU5IEjFSC2n/UDNHz1u2O+2fK/RnTuMPlaz7CJDEei
NIZlzQIICezUtN7QLQJP4LIHX+feeYx13Od7ks5zXL1L8Cxj29sGCcZr6eybHnVWiiGjVwH1LuiZ
t+5SMatnW1Jb0nbxe6rqlHn4AAo0nHro/MFCMkZiHpnO7X+9IpgIVpWsQUdMs1ysTtqJ8dtMns26
Hf1kcf5FenytogpXmPYvnvxKMvXZ/hg3Ns8PrrOexuTq7LJHNclJeR2H7NvuRxgkKA+rvG4JTZZd
gabf3vF/8RtBAAbqqsP3NUSRW7IS3CvtkmJ0dKe2RdJ1HtSrSzAkoJHWam4lmPYr0AtSYy2KNxar
VFf9HMiKqg+q/T8RLtIeYMiEOtnY2Ub7y/XPlXNiVQhgl8u6rTlhE3aYGqbTqinq3outyobqtxcM
3y5xC6FkYrixe39h01izmi9P7uvFrLaCBVyPG1qytAIXxZFmRvLEURn+9igYEsm4hh8DVRt5WyyM
T1OfLoxLHktqs6DbxkJhK/ba5ni29QeiuI0JgNryo1JFB57fM8Fi9hySbuJ1xhFkqC/GJHPxfvII
t7o53FAkMtB0m1ZziWasGj3iLM7DImKb0zLQpuY0YoK7yrZgmWyYHfK+6e3OC15VvQYFbbW/Eop9
ttCfZnwpqTJ6I9r1z0wqrT1r2qHnj0126O9wHydV4tZbQV2kFvi3Os2pxWlO+Hp3ifKjxLMrvy6f
QLw9Skg4RQI8JqRbv0sEmoqNnX8ZYwX0VqSOb8g2fgtVnvLo2weAW8liNvT7lZ4UicXUlStt2oe0
ovUbWG5RcMDC0/ty/bFg27X/ibR15JRwTOR0O4mUtYfhkEMqtsDMvbHVwZ9NxFL67JG3IJdlr1se
HZmVGqGkaUPIJg9/3tUy49RQb0VMEnjvs597fXhdt8xtwx+bLoGqki2XAisivB1Z1c9RPxg/Sbup
lLUdgsRX0vEDj65Xc16Ip1Oit6QzPNMp1fq6jRr8zNJOo+vj87Yshv8asJcGXAV4//Hw4YXBN1UL
OomWd8Oq4eJ3VMHO05NKmOEekUgvvfIE+ytRGMil4KSmtEFpI8ARJ1S30J7YLmts9pBSHW3tRsrc
4XvuaheO54Laik5D45O/Hx4W1V/OiW0JQm9e1/klXCitigniSOI/FrY730V13TNY+cp29k2gmCbr
StPAhVwCu+plrzq8X0+5CP+qqCeeYMuk3oquyHpaahqSdASDli3Rcan9qVWrXzXDCtCGbTVM4CKl
xHCAXRsJHQpqQtEYTgYBxRjrOLjO/rjEXx9OvSMmsNR+pmdLApIArT/8X1d1GHeLrZNLfbbKmCVP
6Y5Vf0L4zRurcYbBLd2jtmuzZxTpSQWPJzUjtCQ2BAGU+MnSvC0cczMGzNFuN7pHJZh3U2CcmO12
AtjkfzSLXQ11njoKlQaSRVqwGRi1YjxrZJiYW1CB+myL1dUZb6NI5um6d5+qQziL+PGkpnTaMgsC
fBzRMNUiGLSPcYcd4fje/s2XwUwSSzHCS4Mlt9Fhu/y2S8q92u/vUpKnDBuJq0gDiCnMEFqn7jBy
SDKZ65kUQ8n+hLSRc7OJQyXIcAsrR/31YBer81KUJcguxi+Wd9V6MhnAkKJp5TecWnkvfEgt27fc
ia/PP8Mc66yCV0r4ZNt90NEpxuao7NBrlrrufFD4IxiUWcq5qVSyO7N1imfrfTtD2Gp8RQILKTvQ
Za2fM91O42cEYfOSglCzk4efc6t6SxxFQXtCuFYPNCqVKbJ4xZpHpNCFBW2ylmtye4nb97xd1vXd
ZeyXIrckfKkvjf9mADS4UB38mgU+aGYB0srfxCNm37VjaQPT2+1Z8ka1xEzeIkgzVA/MbfREwXjm
8jTLS5f9y+Psef1d/fz2Ozw1gQkp4xjps7m//ZqQBW3qr0VVVw2qxrPpR3+lydEwXMlVO4TaSeU4
zsxlO6mkgGffa1SpcDieDH36Ac0J8tV+ha8VRADzdBtqICpPr97PtygXaKkfZC2cql8s19N6zzTI
JOQRj1lfjtFGrvTCjS/dtHLx/IL8sSue8eE1mMEShnSkIazbYDNnCuq0yO/LT6a9oW/aeo2D5C9P
E79y3GpvacOh/l7bd/F2abOWs1Wg/IBiltSNLmpfTSePs9VtIl5zKMHGWrhSZJZnWlG19slJwFZc
yrn0UfHjSAHrncRZzGKdptv5D7szyuaZgpcO1y6Bs2W/OavevsDl5M0x3dybUI9zz31/lTBUx4Vp
Pe/B+bRtg65+HgCikfX272d4u/h2FAooxeFhyTsjmLBG2RBwGElZiKxUGK+XCi8eT/ACYI4T/FQg
cvSaciSBNlChSS7Ub92NKDX585O6t8pa1yGN1TwkjR82iXm1ZggFgGubYmJlzPpavplAYbHvGZsd
F7mfDdp8BatEIPMk5cQTsh1SBYI3BS/nIX86uHEQwlEHb42lzeDXZ+g2GR3Zs3HTIUm8GQqxIfvH
RMfNQquRh8fDbS5Mzk7/DKRGFj4+FNlCVuVHO5J9mQ93TxNU9ZfePVpAayWAu94BRc7GpO+oLzSL
mu4gwrk7KlFj4mz5PszYoK4sIMc7k/ofdH3OLNPxFTEfi8jBWfpDDYB0w/lTTXl2hGHYJhIwlMM2
Mi35G8aN9mQezaMVE8s2UYbyQbDU0RQ0r4m5cqu1xdFSKuZVkXd1kgy0Wh8D4apMpF/cxXJ9D6c3
rIkr09KEvAACr8s0j4THEdcp5oTzlVFhPDP4vzqmeUjtFIXgfDoNu6YOBWyfnTaFEFrFILzjnbCa
6ep3gl6z4babjQC+V0aZFcc591YZLg9zWvXs+obf9t3rKxu0YMdZpYeC/hktb1+3innowKhOVMka
gF0anCGk723K+BjpuKBRl9eWx7b7ILd/oneCQAdHnpeLwbroHYQ1h8voMl2ZCDi6trIUqCF7xuON
9nd7yn20TPGL+fJayqJ7bwMW2pni4iQ7loHDSUnbMJgBpTDwscBBnTZjj6L8CN4f4dAJQAq/X+lZ
2S8CWQrlTH9uFLjp0N5OZ7ryZWUMor6CzaZ/fzJSoHhJP81lKGZJf1HGYBCmNm/XzSjPbbRjk4d1
zBgEMPPF55+soDglN1yo2QboRtEdZbkUOYyFsW0bN8nnCgyrKCerACU25Qc1g8hX5jKjxyOrAxj1
/VsxwcUwmbraE8i8o9T+VZiL2NpDpM1pXKC5FQcrPhI7Gu6UFABuviSE485TnZkNOajpEPiXW9ux
9Zh4FVyt/gDxvZ5IMF93TohcSYplj9eoK8sAz6PSzBtcIblb3hpe/MozQp1afL+jWTPxawB2aX61
pUHyIIIhJyU3T/+ehOIQxKlpMu/r1WAZP7WN3XVXo1KB4Ks06MDiOnf/AxuHfaq85ucXK01To2w7
R59N0MfCKsAw3pgvGh8DEUO+ZguOj1cWnhb9UxDMP49aYn/wvGvFuZVh+4baq9khtR6G8xWTQviW
lAbjdXkOdA3QIDGT55QewjyOgByKlymmoEUSHbEcQGJYQE7//TKquV/TrjLlPBK5sbd7yLcnF4Fp
P21vTieyE1ytzQI4Geg2rdwXdLUcKBs2bRetSCl4pvSDZrHjdAyoobcE9uViqdWsU3Ty13pNDkHU
ET46XeFdFKDWhC+Va49FNrcc8MkQcEN+Ku7t4wFSWnCiriYeKBa4BvSQ7NGFIlZmZn89AM/eYZvB
z/0/AliYeqPYb4fUUil+ldJxCWcePjUeSQTrp1HjIbTlHlBsTB/bOq1W8mysBB9vruOCpOmaF73Q
OoR56ACu+BqiVq12sOEtMyIByl35b3zfRbNnKbpg97fssIwTkw+LuVyR+wY0UYKrL2+jHSytunzm
Utjj2YiYYyNYL3Xc34qs+qPtkgqmBt4lgTO24q/Nsh8BRLidxDKnjvVy3oKxKFms+mYgW+36rNGT
UkwWfXP/G9V6e8+gmMOC8P9Fzl4C904CzJ7YB2EUJlqY8F6mzUJcccrOFobnhF1e/agQw6ymVFf5
yL/HbX/FWF56NTuSGfDbWV18sm58o5995Lvy+SEOXeQZyGzTM+29ZqlX0/60wOxxRcgetQLF6d7A
DE+pNy1PYz0O6QbtknR89CMLn9sTthHnIYcqI03OKnD6lRQbJ0RWwRTOLLJdIUANqBwszSO2AtuE
Lj6PRhmIAwxh18LeDLi6fL4/iXYyGzfE9C/oOe2Zhfg/yCa/+3YvMMhRPByy+3gY7hzyBVKVa9Yw
By4TYSSodh44SB9mDsQNZ7PnXbbHwe5XUyn6NTy8RUZ/hHYv4my7XRMQnBp1AutaewMiqpZFBJdP
4RDGv5gDAJAsrtEnb5ZVTuO4X60KS0Hfnxov7zBOo2vOuekWM6vAGjUCNfQFXBV00BdSoKCyr1gN
TDwTx6GRr/wgJGkwKsIxzqyx9VeILPGZcc2C9iweXb4TXuBzO3rIt9R9tD9MLHjaP0UGnqoFpx2I
SMUPLCeIIqSh2ZgY82UQe6q+l0zvdSGEFd7In8mWCHpL9UFQaZu71ejwUrnmU5zFkfj1qh0NsfsQ
aFwcdZRRittGk69GgxKtwrhUNx2sRz6Fv+HKSA805bwHTele1T9ykyJdfIUVRcN625VZn4g9ia6D
7ZOaKJW3uQktrrXeuMUWtGTK2baGwC8PDDGbRmjWtPhGfW1daW6QfdkC5SbgC9C9vBpnumwpazNL
64hVVtyF3ObZ6tROXLsoG24BdTpJXd9yq6lfV3W438sJlJYeTOUEaNXzDUwix2Q7KgNEIPsiBrgP
05okAkUE9e/m8zyOxYz+W2c4k5chKbQeTIMRCamLUhVIX7svq+1lo52H0MfBG8Tk5rSncmmkYjas
VAYpUcUwDFUx2OEpRfDrMjynpZ44gRrcaDebKgxC40ezYrVXgHhh25bAdyvutth5qBBrNSW8w0j1
Js2mW5wLUkgoh+re3CXChlsFmAA3JB9oV09jT50Yo0E1NV5KgQq+PAwzN/nOh2Q6SSvRNcV4rWRC
aQayy/qAMWrot24+Gfem7/As1iHUEJ8StocZ5lvX3SxaWA8EtsokiokEK07Ww4K/DHUdcDtDfIDw
dPBk8eDJoJ4hOmvL743SOlu/AH9Ntj3uAJJhqOTUmRcUJ+bETIRq9+f/yyxuvGve2SK7K8VvMcqV
+P7G10AYsV2Bs1IFHriefAG61D0aQWrSG24veS9dMA5tp2wMaTrNoO2ldZcor4oyVbu8/Q71eGaX
HESsB/xw30eQ0cktmROpLgVJoLqOns+/6fccCcmL/jzWC71aCi3KiWSwkbeEIFqSq9+vPOi0QeFo
azi4hf+Q7Qs5TOZ3LEj4HCzol5YliUNjoLaLIWFjgVyyk8xmBsk73ppMrRhzzKuhfKX5mnArjIg0
BSUtD77kbEOggKeiPDIzxDR5SlkeuSNZymvDNLotDKll/RHAdTbMg/vLOy6EbTf6cq746+RcC8gt
Tqh/kWL9qBAq4m2tMbF6D2ULzAIGslMbc/eFQoD7mn7Z5xujfSeuje6yid/VvJf6Ja1AT/Wwkc77
Hwh3W7K/b2zRLjjLm0k6q2n2DjiDsdajNNWRcAVxweW7CWolVkYeors2JcL5jS/uRcWraWCdSaQo
lH945fyXQTHujIePtLfk/r/ZitvCri+bLULMRQIf18B/mDT9NxYXGsjtSU/Z76sPYBbik89qQGgq
tKYZbq3EbRP8wigVK6BHf0vr9BJc+5qMbBgKxlRvNDyx0MnV1OyaFNe91Z8BBWfRnzP4RlOgtqy7
8nLEV0yZzpfYgswsDe/DnCrUav4vFPsXiBoFnKOJRhcfip3BRe3bTXwbBJeYhSg983MZD5AK1fnO
5DuMkoBAomaZlPXGAr/9sGjQ1PFiumjRulaeGE47/NSj2n+pUWQW4wxF6Wkd29WvqhGHfyHNi0c4
Wdt07APY+vKdCYrdlttvIkdFhcjrm5gVBEkjcTLcPUCQ8WZMxl7pzZywE5a5+VzBEFRaLXHKESdN
2tJNPUTPu3b2Vnn+kNVQvIO7zkT/DLqmrKJwJMzz0wBDB16CnWI58qEo9w+KySjdfSQaxePZyCj7
ifIRTr1WHB78rf75oYEWkOY7j2T/WoTYdtDT9a0sdt1AWdB6knKWQoP3+kGiKNlGtPvRn2jg+1Sy
FbdpySN/Edsr9fjIqh+4VuVa3NZGijmyuLLBHu8jpzNc1TM51UYvTZxoHXbq3ecurD39ZRmDnFxd
4pVvi2tjeMODJxB45cJTMBCIJwpzwBS+p0gqL8wwjAX5yN1iX5TZFgjC6lsznJ9OMcApj/o2qg4+
NVbSglfVvsK9J7Os63vT6V9ucq3PIkSVsPifV1fm8Zxhperl5ufIZwYOOhJwTrrjvkfaIf9BkSgg
17A1OGJ4EmAQXLZDKCFCLJqVuRC29YnQ56hJmVIGmTiScOlzirmNNmJPLOiZWJ0bFJeG0vnke/QJ
j5KvM7YbvgKe8NFNFsqd7maHWAvyJd0E/FhkMBTZmFmwVgejSK1DIDCtu31yPfJyT0eFEjoZfK/z
pxD3BpAMcOYH04lOlHk4wFTqyTeVsDKaYK6HIqpP4t7hrg2bk59mEmn4ea5JbO4H/0ZLgVGup5EL
D6KAb9MUkXG/r2/jazXUP916D+T9v+JkGiE1ZPeBq/t1dat9DGu6t80/Gcxu9elc7v2Jkch+sjwU
KH2Dmk0PlRPt4wKb3CBBbzC5hzmi0UnO77dT0mwQndDC2EWwaJUCZZ6xK1CDP/XHzWCfsWykFtLo
+kIajR9g+kGYN9E+O8fKAvl6VnL8/5iQwC7ah+z0T2/sDP3Erm1j6qjN/Ir2qB33z5mJ+q4CacX5
V6Wn36kY006U53qFsyaKTas/tBrWT7hPSwVqR0Y0glBG0qM0uIsCAs6/LGgz7RNWVHOOvwX0kDAY
Tp4ztr28EHbUycoB+dqn32X5HogOSeOepjOZaG25Lk43NRh9kv+3NG0yaqkJUytMh0B10jNAeCBv
8GLXVhbdaf4YPUs8gnZz1ElwW7Tpc5qVo9cHn/9H5k0BK7aRYcUjvqNPqk+Y3PxlsJkrb7cRkrrS
POTavaHRuqTHMf152yeybLbVLonMUuVaDcaW6ymKEWggcuoH10ZOOWyjUEMF/T5fFkyNaOtQVotI
1tcElIjjIEfcqCdISOw7+SbJ10VlEhUXbEI5BlrSbtvhf5fu9Qn0IrfeXfFVWRpukpAG/+NVO26O
ddr5/44D76QIFSyu+2fEFeL2wd8Gm00flaZ6PuO5Ta63A3dwtLAOKf91hNzVVFx4Fe33hutCgXWq
fnBmg+SVBWHR4gy7QWir3CIrjk9xVtg/z2AkDBZBRBH6l8fDzF987gqY+geoau7dkq2/SEXG/8As
lwi9HSVDhRocz/jzmg+8gZufGzLM06JLg3jvHwtEugeElJ8j1kZwmZGJINynxeXaYyBFPKYRjMZK
udtmdAggrfM6Y81jkp8HHFVpd7LAZ5cWp3AvPTXeISkMTl1J3vGnsP50kfU3bgtwkXN6HLrIl5Fy
dcTXlZ4vuj68WR1G2a8q9hH5JKg5mwW06WAvhqpSDp1FM/wtd7jb5wUfax4CvjjV4l2+tZIka/T7
fK9talrsjwO1gpufd3tg98CDENgskvcmpSRWW+l7Vg5PuOss2kB8520HrNIma1Y8GgBf4KutY504
z/MuzPVMBWzuqoe+GESwGJtS9JaXsMX+OVRjREHOI3UlQHXhlwHYfXjAxmn+uelPGMuMOHbymo5Z
QFNiGn/us13Tugw3rgMirhv5AukCCv6H5VCL8AwyY/Lz0TWXqeeYk5SNi2Ib2H8oAE7cMMlqi2Qp
ATSNmH3AAlkkgkLMUr+KSCw2DhpJIYC4WxSJVcKrwOoEagWGl0PsXMiazTES6PkASE8dKWSNL23T
EOgt/er9QUKtaPZ93j93oC5pBCKj1UPKjMZFWOw+MtyrBImz2VYIJZh5dpEc1lLPtzx+hrIb6mb2
mMhRxzesCDzh3AjlbqSXEU9EZ1vUB8vCO5AhyvjyyEMiGjOAwq2mfL4soTq2urDqvNKZOYvNzG7T
0sp1m+8jWwIYZxbMNa9HAuFzYqlCS71TUlaSrErHcF2Ofr+sRECuJgWbhlGVZxjq5HjNNG9rSd6p
WOXdyepHH+czsoFFVkktotadyFw6flGPMlIv4KnC8p9x2PmlZnTGnvll0wczWNZs1mAa3fNBBpbn
yYqyFyCh7Eru5pkXp/AHDy3na3FxEl/i9asHLhE6MZAI7K2cUt8h6PSbA81mm7aC0QN8opH7/TCS
vpT33IrlwGF0fhiYLNstCxjnGenYVOrxaSSfoyTiSneGrcSH0+qRf/dSZAxVX/eKS9OHUD8PEB4i
3HLp78lThssvDFWy0jaPR0t/3sWndDS+D7X9VDNm/+0R6E7cbM3+SiejToQgTxpGjKVFZKErExV5
MRdZLKtu3duGPnskKLLfp7sCQ5DYh7kNschATJYZZn5OjJe7qmZAlJTzzNRoDyWm9cd1fm9JWUMT
bMZc5s+/+fHD8uAK1uC6fDOVYSXx4/KLyGOMgKEE5BQjORhWIfzvbSQk/6V7w6qSEOC3Lc3yV2De
wuhmoTRNRr6T9M4kPOLujjTzlEHPeSSaHngANKkm9SDI3Gp/hYepCtnIcLC9bZ7B7a3LGyYVzclE
kyX2SZDSk155Pm+lfdQGcKow++tSPlgcs0hm1BNyHRnjd4QY4khJTmED3o4jOURZM2LkbGXWckPy
BdT/CqEgmJbZJQ9a9LSk43pPmPhh6dVRhdOReY2j+lfBHqSQZtM78ioKMZ5+v71oEEciopPnWr3U
l/tuA0cz39OTO7fdluhOhyF7YBZRZAGy7VjtaEJTV93/Reww9K9gpudNzptkIwv4DOtd/a5mqp0x
4UndGU4Y+9CxZBXA+5xioMiiA6ccjC/OMOkDxY1fOFKjkwAncU8eVmDPybNFUmdljGUN+KP+Y7MG
Z0Nmpq6pqci50Pf/Ahg3ReB/y/X8f16GlG0ve5DUX93VlRjWc1cG2yj+YKsmdo7cpc0EMSNnun4g
fKVJ5MwMkHvHeh5wFGnWFaBqX+W5rah/5yWKTAswi5uey013r1zFNktZ3LsHII2sx7WPcq7qerTO
Ti28Kdeh8G8OjcY/KrSBS6Zy7qqmFqcpFFK0V+l/Kd/od9y2+MuR0faAbZESS1yjKdzxjvB8uSxf
fwiVaPw2FVcJlb6fle9kFlTkv3ncFts36h5JfpZFrLxSd8N05y+KY/pM9VVo1wdvu8HvE7kpZLAR
CSLJiGuK/zFGC0yPrPMaPMPhm+W794EYFGzPObSko4llBL7PEpHX//kiZmDJ2vcnGdaE1FX5pSvi
Ix1dhRREQfrGVP9g8Qd9eOyfkU1JAzE1mq6BbCd2JSQrmDx0BT5kclSYPPg1IPPjVJ8ieyncjNtl
5FpOP5Z+gbDe8yNLFjm5hDiJB16A0dnaNi/C9Q84hIzJMV6nIvyNEvCu6kAQd+9U1ykymKjemy/X
9g6UuM9fSwEx0y65kumj+c/K451aLKLE9gIgVydXj8IOsTpXZxl78IHhoycewziRmTkcHv9CGWqp
eKjNEdws5MQBhhlnyGoGj3QKcc7PXYC0XRHz2QnypzCK/nijeHxmg5suIiN13gFcMdBR0+AFf6kC
A917nEV6yLowHEQSwP++BQcFL+UHbTdnnyUbK7FhKqt2EeYc+bmua8d6EW+SR+QOGGIZNo8auP0f
vmqGM3Ztzx89u/tjHYEGwN0w+RwwrEOdp+Uzk8occPsTNU0QHuGSA3D0YCP0gipmX2nVohKqIl4S
+6LOTwdTM8s1zGGEE7LTGOfgv6+q04bP29ns9MFIFArR0nC7nPHrcWX64Wf4NQ4o+sasm+gzoQZN
QhkXYwNCBGgTRtvV6Sfuj8p6/sJxY6Wk3WoncVkBQSHSAE27VPZYB7ncrUROLPComzJYTnRuW6Ns
91ffYi9Ww3/uS9FI+r/YAvhAOfveKdzCOf8wC4yD8qLNXGCGW80ZaVZ1dOZlgX6wYWjXwe0c4vN3
MaR5h+41w5iW8vSc8xRmIrEFNb+yOPMW5zjLj9mGowR+EUshGU+EYZ4PYDAFlYZhjhMrwh0tzHHp
CWC8aTP1RdoRK4dEM2FAnbS9TjHC3PhcvszENBXBMKJ/IfepJZeFYmRN85h65V/OP7yWaZpABr2u
6a5ATGLcga6lBvl0X5QL1kqLwndSfnapcpMGAtDPVyvE8nOq99c/R6rzwXYNjHvHBOaYUQhqlJzW
yoNL4vjD3qBBrjVUbVLq09OvUuhshl8+dZq4/mIetXcR9XFsYLhisXhGyVDAy1V97LflO74PfdxT
cp/yMNkOn83nZs0+2D7GE273BLxvjih1f8/o82l9svHf7KR8FCZt8DGdOiAqT3I1MHLcVAiPMRkL
bki/bZTDD6zWwpY5KHqfabWfulPTy3FfBJaqiUPUGoMNAPyDinF6DxhXvaNd3X3HSLgoG2X4pFnM
VVtsJDi76CacF15epdXWfHR7rSYcql57x2N4+/8weyBHJdi//UUJIrEFovcgBGBPZMFcs+Ef2vtj
BCjRdoY3dKxWvST5OuIUOBGJcu6D/JDKFwCOP6gkiLCq/zDrYs/3xA/w8gS1QU9uWSVKRtANbDAP
HfoGX9bn8ifEGV2+SKZkdLFmdzq7i4Xa6Rx3lhuN9qkZDiBCHIHrl67lN95b4qah8p7ijgwboN0/
YdueyUh5kHvD46X00AC3tWGMpezoGHzBPQ1BdHKQh3NM3Clcaz+wmFZ0Qmo5Coz3O/sQTMRILR/p
csCtVH3gXHGRdlBxBvo3t6TQlGXi1wnwrnrmROAR6dfnqkOWgjCuSLHSMsaETh0t8/QH3Wc7esHm
YgYQqoUHCaGtU/Fls2vte03ZJ53SmUnC9hBweJEDs0QcZran8e1YeFGZ19m2Y4CZ70wPo523IGpN
aXOY5COxreusBPAMb0l4turbcZILlZqri4JpDDCGyq2WKVcCYSy/0XfPXMk8a/Byb6492nfSqchf
kSZwA07o7Y2HdENsDraAA6FZIcaUt6jzvDiVw7cgEyovaq5SNY5ipr9ueGuvX0xSgviISB8QBmhX
6xUwHbPK0eK8Xw7oRYELFOK04YHAQ/kyCbfH82Y3P2qH/4pFfsDyACflG6ob4y3OwxkXffBIzlLK
XEKirmdijy3DZZI+ZrfobJ7hqTeyyns4hySCbvIZEBXN7UffR8LMSgIAikeA0oFCA+M2fZT6RIb8
ttjyUwI4kTYqNcdNNExjogeAzUJSgZ9xqsPMREM6d5/ZXCwXh7FXbSfy5UWUoWMLb4NZszBCeR3M
kLZr6rM/z4UozXPDxYwCcYYmjGsACA6JD51O2JkMxIQfuiYlSAOc18i70QzYK3NgxSauV5p24zNU
j5t7dKshUE3L1k8i4OWmjHbHwkJbnRZ6td6j4+OHintiKqRdx2uhAfOaHE5dL7zYSQKmVn2pOWtq
6/V+9NfqeMb3rDbKoNxGZm2XhlAfmoIy6hL4M9ORBBTUcFIzAjmeptjmktlaInn4uSNKChMyp4Ee
Ep5pYXze9TSacThcqSxFdKos92CYk7BzLCwan2npTDFWyHopovRTLuMhe6a7fJWRm/1ajzK2Qho3
4g+35rHAxJgGSgUOedodaJSrBGKSZAszbU4Me4cytN7Kx2BZs2K+p6dpDnSmSQm8iRULmPWr5Fom
MdUfUbCGX6yqTe/QMLd+0JUT8f62vS0S81+DAmp/F2rHCtoPSHT6+LKttN4PrQ9yFsMjohYQqcfo
+ZcN4Kw+X9PwSMtCpTxL/B0EyDlcKdT4Bx+diUeQh6Zah2W7O6to/lBW5dTwWI1MD7ctrzIikLEQ
wtefdsIweDFm44sXqdOOWe00vwpFnw63rlK880Ht9fmP4xvRVHaAjGKE0P7NqSC8Wl19MtQ1FayX
kY58e5FKIgeWweVXbAipGJEZQUDf76hoQ6QnmjRT1i0Wp5CFxZkaLHLUJPaBO86efpYF+smdXRw7
bTnrEbi8jEFic8UeN3pCXS2qSvdj4rNScEIDNynAtWug0kFt2NQlFAjOQcoFBG1dDnM25NKB+qcX
BTb9WGwglDWBl3Bj9CqUpEVWqewW6wwRy8Em1dSsdIbF3gm71jNGvJkGLQOhma/0sZ9D9WZ+l+Bz
q06mTbawHP7Irja5gzze+HFdkAlkFpePVz+KurVG8TgBbBRpCuEfojQ6+fPFNRinVnRMdJmesZ+u
EpPJBTcTKq9p1xdM7G7umCXoEAWmymPU2iWKbDjXKigiuHRnMGm/DSRgsMMFa7cnx6us0dyw1kZ2
S4KljVQ/86u1lGf87pm5zfrQWFmKDcCwtITJJ+yE2kT/kaXp8ybZ2xPMLWvEXw9W3HdUIrdgWYzC
ds/xsKG+r1hxNSkb2DVhoZnKeoXAIhQP3CPfPYYIk+XlSKgrye6xTRAT1UZexpaFS4Ep8TOsUo7N
n1fpIHXY77NmXWe9XxK7CHENVsi37pUMStAk0ypCHmvkXOnOruZ/DBQm2ZhVUN6vRDhKlEUaa/Uf
LI2UMp8Hw2pFMlaVWjY4tARuUmkUzD5AiwucdHZ/250BuxFd//rYVgUDwRV2xihDlnVgTuMlsRMB
/60imKrECv3hzilyDParM9/UP/4TXfyaG2oFOMuLNQm+qbMt1uP9XGNLCYPKEgZiCLCsQfUp0KML
8Lua5b4kvUEliVp5pZ9cOzGilzn6wSDdYxIyX5USQVCHFYCMf4gwCofAmDrGrpL8nATYlf2pKhTd
hQrYxrXuhP8eI6JGRNadmp7p2i4+S3vHf+buACBcNpgzYkTHZxaQ/tM0ZU387dBRr7NgLsxmMEfA
c1czBSot/cVSOHz4ycG4wQ0qEJnosPOZpylkSa7RL0STMCva0OfsHEPNmisj7E6RLPTxvIm8OKRA
RzqBz0irqIsJzRasJj095KCMKs+xlo8+avIF0PX4p3TvPKfzwVpnotwzuSgDdvOHkPiVdhRG7Ib3
vpVMa34X0gpjPdsUV4BczRRZMuZPAU/pfSYLlYbo1kDsqoZ1kG30WwJd7Tuzg7pbFWI5obA3taHi
ePTgdoF2klB8B5eEOCEqQ1/kB0Z+0KeUASwYtfkoR/H/ePpbGiBQgfO+T7ElQnFsDmCRtp9yceRz
mFA5BbKFcmaK5cSKgyzdJVqYjhxfFdbAUmer8DgQ1h0SKpZ1hb+d3DxKQNNnJIzfpo8OmNo010GK
/HHFSfrvD7/6u5t80Y4zN4yR93OK9SkOlqU8rabvuLh+MMUavzQ9Y2ZJ48Tz2yQXnQrjMaW9dSlA
FiYnlrhiDNKvdd2SjKRCrRvIQM02mTnT5YvY/6ByGdCgDQA1SBnZpUBOC+NOe/OuuOZzESsTvso3
kJH/Lsb+JHEOztslqlXaBaSMuQK6NiLyOLBRU+1WIQKqIfs6yVf6FBtc0U7ryn6NBeJ42y5A+7oj
pZB7ZL18RlMGinlbhXkbIbJR3pmmd/Mjhh2fDeMECwWyze/8TkOEYEf93uegHxIkqPCmKPmIQBlh
2XfnuLlTXNvIyysTEEjK17xamqxTHueOC8XbAsCz04UfdsrDd7rMQq6/DN5QSBrbBRV+51ZjNgYc
z6v/CtSQOSeu+Pulwy2DXR9eUptCwlP7Awc4oIgst3UBeddBXTqb8hFVPjbBD+xJG1r8YvaXZQ3b
jNH8YzdJaKGCvbLoGylPTadXNrUWgRHPgg5DJlvWoooUQnWbh2bJBZPyPGP91jWRSQFac3woK/8w
9Xx2A7zYvApP38UEtXeLuSnLQ8WS1C1o2Dy6HxDzCN1e2jzZDAxchmpA5De7Lf2AjiyI4U05MLjf
5nqm+P9lPnyJc0DFISLDp/gN7wyVT8uTxl4I/DXUFPRExtsd6GEr3hdPTBgh+XaUjpUPe9gBe5Zq
yHytwwU2VLQ4Sk63AjUwQZlcwTBNIrzzV8NKJH65zfH+HWa7h8mfA8WVHRhxciImT/tkX68wjfKs
MC/LepJRyNVFWIDVP2OEkRar57lQBFaeuT4CbI8tBv5iDJ79KZRxxRbfE1ueAhbX9Dq0HLwiHQRI
4KVwJaxejacsaJqSpkSfrnY/SDs4jpokEQma+LZoDBeFp0/kyhFtC4UZxojBXr1hFzL11EueOTMx
NQlEPdesCjTPDhE+cwVzFpLvce0C/QLP4nHfMeElU2U7fL/cXf4lGKh/DQ8xAKhY0Z1kiFB/1nzW
hbiEGqL2nAzDEFK+8FfaAjvjKfRKTDQLk1CSxt8f9OvCs443aRdKlZTZbXb55HWimdpjXpLEa07a
yEsLZarkMiemWFXOzPF3xh5iKU9pZ1DSeFjUAuIID2f1TqUkdzmJL6Lj6DYhpT02izLf7NkO9t6b
4PMNcpiRjlK1qmJkW182Qtq1Av0WAeM8XY9cxWilCdtn9Nlgp7sGXC+tzkw/aZbGyiJViI+qPpm/
+iWuq/sOVlxH7MfWgMd6DkVbre6f2/tshPKeT6IHtuOwnWKR3bZ8/Vhf2A7DKKSThNJ/WHXfYMID
fp3Zrk+RoG8lP1MTEHR2uVWjCXcZ58IA0jlWGfIlYI4xRXWi31gBl+5oNZipS1PuVekgwoYQBH7K
aR8GhCagYlAF9yNrSAnacweVuoo723qJ8p07lGpuha6rCJxOiDv1E383e/yWQrZ0gdD+og5GMyqP
joFc7oxRBbyzEMV08cAWPnJ4e8fcj896YqUXkf1QYiM/lYWtxyI7VUYLyz72iPyrVN2+67sJmrcB
QXAa/pI9Xqmr4FHDZl/IpsMuQsH97TF/ozagnDDM1p9a8GAwHs7LiKqgbgcmfVmEUAEkeieb/gcT
cbBfyX4mB9PlNO+EmlLKgNm6RFwnX6MCWeRzu9GjOKnHuHB6E2n3nJzF8zZ1+Pp1VGB7xQ9Qt+oo
bKl5itkMtBa3z969Bq9xFTb7Po1qlhz46KrbvTPvbSpN4Re+Ubi3uWV76rsHokT9aJGFR5wX2NlP
cJSFwE9+MK+JSzQq/heBFwXbKMR22td/tohpLFe2meuRa4ezTqAavk8fnAU2W8qeQXuTfVdazWBZ
6EQ6tkcuXn/JmjuWUXDZSd1CF4gDF3XZzuNVG6HL6aHSZn2YaRoHReySvSMLEx3ibQo5zsGod5TB
1ClKzwXm3gkm3kPwXBBNoSFhhxpOuHLLQY+aSMb1w1KPovv/26Y9vISLERiiYtecbUDs0kbKo1R1
hEZQ5I/wMQavcouljpb2bCg1m1Rn/Ngn5PHzZGgOSwVOU9b5me5YDA2uJzal1P4Rn9yNQWiq+4+O
GW6PyFFeEGSMVo1nKAXOyTRG+AGzMan6T2QzcIf5tSW8y2N2/jeokAd6m5O++xYUBAf1ytS2qVLv
jIkkwyMQzu2c6y+vCJe9rQKal4RdTDvF8SJuyVb1cPGn1efs4yR67avdZNDbFu8h0iKIQB8mfKWa
duXNzE7txVOaoQnkY9L5F5KXp9IZjolfVT6VeYgdMLgVgW4mhBQq/2MsgZFgLVdtMrZTKuCiwUvo
aXZZXOp7zrUj+ua1mRKq7R95FCNP77NuzswGP6nECEZeI/jkJikBoZZtbsTY4GnadwHUxsLepmS6
ZMTltg2AYTRDIaviGL75+dZaxDO8RaTMulHuxi9eTYg+XrEdVUwj2OeFzkDKrWHLjWjn35GQedTe
OFMcVCSQVfe92kxQlU38NISRDH/aiCKbi8uzQYEvGnZXFhvpRDhgilM+0JfQyOnWPXs3I5kKX/BG
b9UgMkGwBXPxLc1IFCkfAtDNPcUsi7Hyf9IY/EzBjLXy67djds5wI/gW5QBk1kCr/0M3LDczzeya
1GR6WEE3g3oB0iu0NGlvWACAYMpwUjxO8kF/r4cFPZp6f3CcmjHCsIWkXNux0d4ytSCSoTdtJNIV
qETm8C9mRxk0EB7su3woZSlI4Sq7sCQ83XSlBwfnx1NZfDR72H/uhpI/IynSaK9fZxZ87Pv02bn+
+SDg4uFLj6pdZ//Grptzn9XC8JWkKNLaAnxpj9NE0SOQWNpYxc0vJAXM/2l7aJbnMxFeNNJLkH3G
jHwk4SukaBE8A1nlRcSWFx91X28hGD8uObEQhpYk5QZSYICyje547XLUQ3nipKVpSadkyelEIdc4
dRHSYqFxonfrg+XT0C1135WkTtsRDUqchb5ie9ThC3R1HXZUF1deeIt/Y3x8IW9g1ioiQbRY7oaG
BTvIZrqgiy25szOB5+5B4E2CkdsVAVjjdIchkFI71qMntoOWzw8MJgDszY+OMYBPqxtcaAKnQjqh
COWiQ9m6jCMmwqI2ZTlpVp/n1cJq+4gSRofeahiV9R6+DO2vnEarweWMFx38mhwEzEROyHP+RHS4
mb8O928vXyi8nfcQ66Hv0TYxG0MBJmqbKsyGT2yHX2QttCFN/iN5SJH9ECNAKeSOQpqEQUvIJRWK
VUPDQzhjcZREJVwaY7PuXuI41aRrw1f27NE4flhvnAbUn52PypkQmclSKmGvt8DilhMSDxoqbHSk
7E/oGszMXnzZkE1AEXVhEkCyEHzfxiSZT+LDY4r6YneMqKaYnySRCGCwFfARnNkCqe1M6jkbXhlv
dvBUUJpTcrKTJ/HSnUHIAPOAT/brCKMOdRhZUWm7A3iLHSIhMqY4U+R8Ul7hcH5PMwSMGK7YinvH
WvGuxaOVkwJD83+Vix3QBVySVJVg2fRVu9j8JzruOn9QKImlg4am16y0Z4QPKftTzFfWkN3WPEJQ
ZrYThUKdUx3+y6R61AzjBGKCulONySUVSwibjjPBM76qxygMpl0YGMqByJNjSihuXXJ5fwi0VpD/
/k2hMffnOpSZklwEe9oa4WFXBvq6vFzJry+slJGRLgdPoObnikDEgbytqnmZcg36JBsseWEwalke
k4/Il/V305DQJd6upu7WsQg2xOj/vj7gl0BPxxE+hRDPaY3p9TJ7IQ2btQd84cMfHh2kHWMrfQOl
3ON/iddvMXg/PFCmxk6Ch+1G18k4tYlH388VspERpkhFafbu+tf2bF87wpA7NOIbcamTp48ERsQO
953sQCdLUcTOBsECL3nO0Rz9XJCd9sgnNADJXvx6kixRNiEUo/fAg/QXZQrXmS1FUUdjm4O5iePi
27C2OCreEVL3hoRLVSPRXtqmLR2l71bFceSM0BASKe3qb6wAvDUHhP4b0sh8OdVO4tUtEuXNDfRW
IPxa82+ob+mBYO4DbJtwdijz6LJeMJKVNG4AXdUOXIWlf6XmToNGatkjGGOdnL+EwxZM2Q+ZjReS
280H5qHu/yG0KK6JLWxKJzJ6IISzoH6SUtfBQwzL4YE4AC3B/MMhNa6HXdme8a/zcqELHDBk5OTy
awpUlqti/fe8tDKni0m2SluP4grIyia5+djlE27lCTmFmFra8N3qJ2ub5j5EPZd80V45FcYumX75
acq4yqA/SSR37/ANZH444yTEwi2cYkVZZ+lvqrjfP96mlvyzmMKzqUsrkos0T5nxX0i7p+24jQlD
WPF4kRzZP8EcTEMOTPqb9e8TibcngrDni6bHBvcsIrjSWxQOUhMyW4J4D6HV764em7j7Tw3SioLk
XgdUuUy8+JN61wgyVLgYMmkGls5hYXTWnKwSA/5ScPPpeaF0Bdbpk1KpNXzr1fGr6l5wAeSWqq2O
325Er9kvsXBKbdEZLRjwcllCHWYxiwmhZvpCKGi882kfikqec1fSJWeLAeubJ7l+rHL6LX/1e3JJ
KitLwJ4dSlkpByop5jkTNMHqrj9Cvf63OTbDewEHwUO2YHUcxb+19ksC5kaEkbaljnmdj9ArbRbt
rsrxF1POiGokXeQJ/VXArrI3H/vC92LUxQyDVhFhwf3NBcr7D4ADAPGTwHa3nkX7m6SJCVuIn5Zt
R0ZMJk6D2yKp4dT/AbtPzVJT5+ondTvfToH7u9Q9a/S/WgR/we7vTcDnGFrLX8R45ByVBlrfJZP3
lRbokBbK4OQK655Ejld7Coxi9EyfEHeIgF5HNK+ojcyRreXJD5HAYx2F1Oj4XgB3JBG9K98NDW1p
x9wzThI6EAQOoNFE7t8CZ5MSMDZ2Qv7hry0FKSoQFxRuHERQFxvdTSBpS+trXmzkeEOAqmzalC99
smr78fkNjDylUJRlrOuAc9cSNAfTxtL+MRaLfx1nilWR4FgZTaEg/CEZKcDK5hnUf6StpfhBm8fj
dzJqx/q/qMFJB6cKqtEcv1GTiKzMo4NtUBiMjShM7lp1XJ0FSV97hkDjaWkIF0xVDJYgkZtzaN5G
1jwiWSC/+CECbw09mUjfBobXjkoaKEo0v1jnhCzwhOalVDA/Ba22DFrLa9bC5Tib1cY5uxYPo5pS
VtDBCmankjmd/+wD4JdcwYOgGuBxbTXlAVIP4cB4kF48CYr6elXDTVxVEN7MbcqipjjNhoQtl/Ge
TCHoy+yXg9A531EUDM4LVEn7OL0wTE1KEyTI7HgRbI0DBzp9gl6HHAEEsmgJMwIW7UvYprzDtcQj
ERM8yA9cQ7yqdoP6vDZ2s/Cxx+A3PRkQyqjWkGb8zm3ippHGKUrRiDar8RG5zjeCrz4RNcLCBxvB
B1uLQt36D8rdyEMV73nNgrVBCpg1VYAIaTTEvFaO0QXmsIk659PX6lxTzejw2JHFhHIORfidpdgH
ytqx5iimi2JDIhdogFtk/+HUj60ecj7mRQ+Wfk1utqRZJnMiQSxz//G8KE9nSOg4NgCfrhq34f12
Cyt6Y3IHpfjS1uW4dxwBSJC3V1KH6hAvSFbtq3/abby8nnErUUWCaXJCQbDaMlUbFX1hNXpv2l5W
pTkKA0CLC+sfUAyfxzSromBW67zSYO498VWsWAFTAmV5nGCH32bH+guklczMicbevg9v+aWRxPuV
+crRd7PRUjrcKqoYpO1X82qjIa8BHCt8RvT+owltcS8j2e/P9zXjtBOQBDGS/pBGjzRrM4niPcWD
rAQFLABWcz0QxX+T4K/LCwBxV62bRF3/JCxFVXrXW1MOWpdQVZuNEzv9GIoJfTOHEt4mgmn+N6fF
fxp6BK9E0BmHOTijVan7DIZajiDjbWatp4hxNC9RSL8XLqQdwQ1NzC4LwOrVMLhYtcNsyOCvKgIP
Be9ES2AQynneBYCLmRRFerIbiERDggrg2PI6xip5k5CF4cZL8zLyOM5nY3ZojyeacRjh7kn6liRy
rFelpH4MGhIg7ibXXCanEJLtrs++VMppeDmeLMalZDpBrXwIN86ATMFlrYEEU+Dy8uvXxtqevCkG
wbMrem3fgbPafxciDhxBeft+lZISF/4KF1s14XLsVU9qYYUXEJ9XhLnZRWXkDegIf2yvGfU18y5Z
b1E1qy2XuMVjgzD1EOyBE7JI3DCF7W3ZRPdcbJnEMmZuKbQMmdVmiMmkj4rb+fRDkifa4zPJ7rpu
GIBPA7DtazEu/lLCh8xlyRpCGNmPflo2X3Xxw4JfKldIWLohJRlByc7HQRijztFLB25UyEs0W/Hi
BhzyGyJ4ZrSgsHYDn9nTlqqxMbyO5+8+pdeesdvrO3q9wLrKuyuCgI+sf50nEJ0CBP6AArty2Zhd
ridHVLffZ34X2lj3FrQ4QFenYO+sZhaQvxdo2E5ByGsqwuTWNqzISypDiFiN5FPXiVDJejOlcXcp
depkVefEyCMiDUijZR24YY0pjhr7bePajg8ACgG9kHmtKbfmCK2rQEXfjzALXQmwCwk7mXNT6MuM
dkao5HGDMTxU1L21E1Mg36dLPjgNfjv6TxbkQTWEig/+WR40wXtZeSOfTaeMcqmbJoOYN8B3S3Qp
a00MT8arl3nw9zqT1BZExZiF1L++tpD7qsnd8AaoZBH+NPcIqd2+CPmUZH0FqmyFXv0dP19JYhgg
mm44KW4nIemkYkcRLVn9AbW22yn98PGyn7ASKNuyIxbnfCzPhQlEIk1teE7ggnqWaXweR2MWyk9+
78I5es5jXv3dpaM/nO6POwRkkqVFXoCrmQQvhqF1iyDMj2RLvqHurIjDr4wN0SBwUmNE7xd4PTgh
oRP98Wyil0MhG8jKzMy2Q3DN3qGQrYc09vtxLU3i81Vvj0cEwlLZcj6JsxUI/XQz0xDISAG+jFHr
mF7zcbz/Glb6VlOsTqdQ++HXRKW0De419rJ/cy2ZK70AOngo6W2KF6LB2KeFj5s6IM+LRgKiDLKp
kbL2S9kzkV1FJYJO8U6RGf0ECj1NWpoKKHUzTMDRozb4zZHMIk4Ywwtq/TO0rt/IJmxmmLaMVS8l
wW1a5M7uDoudmzbmcpzV+Y84hX90y6bvN8Vr9sfZgyHW3B5LJ31knrUq8LEsgHrZnru/nj6d5u02
gus0YrmW60Oabfybq4NYg1AgKKi9kJSCcY+9oo34R3uA5bf/V5K2v74Xf6wRMsJj/ajiUysqzGHN
4zdrIpB/zw5txnB1EjAfD8Oh5slUr53+mMjTz5Mi1NiWdKWQF7ji93IPafKXGmOSAGnI4Ea7h2di
NUppSUdB1YC4+NZ1J3x8JumXHj/tj/YS0W6kIC0ihFndNLNasVZN7FgolRXYQOVkKi8YjAf8J6bk
SdOXpVhWBls2M9I1XqcbeCSFkJdDQ8hKDQQV5I2xXAnpj5Y6fUAv1854cny7/Z89+jMkLq1QQlRn
0X+fL26DHzPoO1iRPRa74fQ1i0I1oalCC+LJoVPITtllpXB+6NJAC6kQ3yICdGDuW00ZrEv0PQej
PgiRPkjW2GUl1jmCcYzn1le2h/ND+Ay6t3PLZxasAut/Yq//ph79RpcN+qoh1YCm+xV+DeSCn00y
isEdgKTLM1ZkhsC7KRuqxJCfX09pVHSWPSO3OSiXvO8gXJbBzctsrwBSXSXNfxifPsfbFFvlYS+e
zJoBRxhoiM2MgDVlvcPZ7Tx9RiND/wI/ROCPHeh8CRaUm8N4xvIROq3EZkmwiM5VWE6iKBSPnQOG
JOSxani3gNPGafnaaKGCeXQDrHkUKAl5WUYVBCYCEzM+Et7TPB0eJzk8DKvC7cWTMuQa42wA8y6g
qPt9zURyLlI6ZksV8WIeMsN+/TGUM4H/ZyciCFt4Bi+dkEefIbqQXo8WijOYLNhXnnrZFNTxGLaJ
+MTb8UKsIiBb85SwNLtM4UJ9UOZnEk/T0zElVk1ISP+aam2hJD6uIS2N7KkY47V8I3dCJrknuPQY
OlGocLmscQzBGHwoxsTSVwlMBxGxEp5VvGdvDiRJ4fQsApl5ku/zM2/p+b7z1VcL6G/szad+KhmK
OINdOjbbSHizxqtOg1FHpYN9XM02vZapoj/0ax5pQ4cgChjfX29mAzrpp0HPuJn97s0Gx84G528D
hl1Q8Y9gdqoOOzQAomhlu1sPXA19qDlUnr6hrFbB9TXgMkChp2jkb8mnFAr/hIyowYd3Eo0jtEJF
L0DzKh6uo1SOXgJVtjVYx/R3HuTICpZWxjMpc5T/Ebs081yhIXQa2Ab9IwicI7YE2LdFuXMonc+B
lF7XcunHCFFsINVexLdGrAkGKEvYUpBBV/VDA1s7YMURCdzXNdKU17KkanVsPpponvisqjP34MBj
GgDMB+vJA6AQ5hdUyHhWduh7cfewcHNnNoVUEjW/RkI8Axa62IAsNd7fLV4hW46a5q2fIh11qYc2
tJrMS17wVF+ewWwKSDnP7sqpKT4Q1K4i/MfMtb8o0b5jZDS/tQUlUi33ECTBmMw1h3XWuZA+gmg/
r5U2/fLlzQe84Hnsnr8KlnMyjSoJjv0fUwAX1by6llzjeSjNE42S0jzKcDGhTOuZpRWLn8NM9JG6
M545D2TRahPOPf9d+TCRpwIVmg1ZJ5WfxOCw7RfBKxsN1/LU04EZ8HUN3uPzgzlDakJH1DgYrsnN
iuj5CIKb0OzToj98Xf7qkCL1Rbh1FQyUtp61tkvisExEk+eiqjAk/jnGrNWa8scZQkb11E0h/zdD
AxPxjz6z1b7NcUu/ioOpcM5MSf5o5zjT0R9iwOxaLC7p802eaR6JhakqXJIrndzX0mtYGLCS3G8a
+PRlox7ola1pAhKTBRQw1ZS55lWQiN5dUJL2ajIuibMyQLFe1f8JQDnSfNCZqP3/JVcPp3rwIsBZ
TTl01cym36c8cPFdSraHY4OSCc5Z9pSMluWoQ/s+Bg+YEsQlUbBSgJa0mKxLH+j4WjXbk9YzvG8J
ebaLCnApVmIYjjAXCd0Fo2h2jqsi806qlOWED2QWqL0Z4GXmaZaV3svxETE4o4aCx+lxiqwRWU94
6+YI3E3pPXWWgEMlh1tTLBUJXeGDtqSlCOxPf25kSbzKno08aN1IEKlcui2nDaBqI7UcfGk19Wv0
q9uFfpn237VKK39SJSdRMo4Lffy4nOQQpMP8IZZNnoqr2VKW96unBNuMV50lS+f4Zb+hPXSmLGGh
B9JsR80cSC/y2hTrOApOnGKT8HsMQY/K/nWGJG8h5tKlWmaC1HluvNGPhj7wPHGkU4qdqME8Ijjv
ivmCGD/ytQHFuB7H4RVxJMGNC/DwEKdAU+f6SkK0D2BYdqv45Q8CUNezxA7hqdRFaD7+znXiJmUJ
ZObDYo+6Hr0HAsx+Tgnq3y5JT6kh34ZCWKdW+W7aJAnHh2qgDTXTmuZxSogKEi4ftl1RwZXBFPpb
7GcRNxprtuU6a6QIRTHpVCKpCJVmDBHM16q+9D8kUA/37vAQu7l3XQ2Tb2L9WtJkcGdIZQrDNeEO
e32PzWS/cnnxhoZUxnBalTP0EhrYvU6giWpWPobMFPbQf1lYRAFLWy4RQU6mdAN5eq/cW35eVMfq
8LR4FecCbik3eaH/6GCyZ8I+LTc6t7cQMQL6Imj9tqeGkAJaf01a457ybBF/T3aATu0KPEY8s2H6
CQsaoeBbwjTiVgiseVRJIrfu28Vt3vbajnQORVBR/2S7yQxHV/pQh2FMbbzx45VkCI4tG5rl5FQq
G24q/VVqPa1Cdru6EYNdF9NwUAlr9P0KT3kUCNp7MxVsRzQx5QdBXwLsmwUNqTxq8AcygNU8+6A9
T7h2a0G3iyQSHaqGGczNCRRiTqQ4z6NLqz7wCYn+IWUfMEVm1qTwSo2N/4NLNlgqdZKQ3xPBr8HT
vVmWLFu9F4Zw39sQIw4pecHhy6F1hZvnHm215yUkbEVVwAeJuI8XDxDD8WfGTI9aq+ym42hQNKCT
WRuLSB++05+YS1KgypDtToqME04TR/8bCOHFVdArWrhNYQZDMkPkjW1aU9a/QmSbe1eWlp5RZLdM
XCCVJG2Si/2Z5Ulh9MtIroMRm2Vpr4H/vh+RMaF9kmZ82F/ZHBPaRlIV0Y6RAJGLO79VbNipqo4p
u9hkJh1tIEnzI8k08r0lC7z3WX+5CWwnNzAVURjE7wgj/2YyjijEMD+WU+a8WCuG5Mg37EVbJvKj
FGgq3OZNVqhNE+g4vt+fUOm2RxPFfl0nPGtUmhXwojzfm29y1ZTy8ZDD6X1mJjov+P0Hvyns7MTA
ks1chfP1CJ1qqRa0QQeMgx7S8cGuWX6vw66FcI/fsII/Y853IbNiE4ElkrkoDhOFYYDPcVc7o9qX
yp6KaSf/CQyW8iM8v3NgRG/QKBrLbLGoeooQW7//V38r8UowEqiexXEU0s3pJfFl9EvdHHDvb+4Q
asH+ZQfEqdyuvTbQyj29rnEb2CT+yg/Eew/BPruwddkCfbQ2Nd0zwoPdTKMODjZVfDboS53d2Dt+
eRFPGDb7BJt7/cV8iPQlgm+DaCCf4+cP/ncOeEySN87PnB0ExQc8g8rUhJk4UOs5NOcNTdsmXwQZ
vLvdqVZM7KELxyCVABdD09iqABsQzM+5rc1xcKe6hc4hIvaq+EI67H0YRaqYVYNO6YLruJO3sS2g
/SG4a+IbYYO8RvtlLBMZ/cLWn/I8UfpGNTWxDA7yUeG8o0GSynoCdBdJoqCgBATXbuA5/N/W0bc1
VF8D9q1k/jEGxjasCdjSUKs6x/QSOoKNl6FBBv4m/fIw1+BZpYzQ6r3OvBK79hHZK6S0Xux1hHcJ
T9yh8g8ik6B1xhTVs+uxPQCEJcwaFdyDbJ/vLmXBSvuHa+TP3/z8N+J3cpoNjg4UuAQEKCdWwUSH
fvpjwTdsUpc1VyE25mvEPZ83p76xdNpEopzZNARQEWCtAmjhC6Itp/E3BH1Q9LeEFWuSWRR6da2Q
vnhMUK1cGaBfIRnwQKyrhEG2KYHfD1fqMIUscVAOA84ua+smnxejml3O0Ic9nH5P3f6XnqmYkZYT
p0Chf2YyQ0hnuW3C08FPqm7VsHI0xqgUcuo2HHiRQ9KDepyRIfkTYiKU/e9un2Ig06SmLMbfGU2+
rh/L+qxsFm9bJJvplqzu02k2D/EovrOYTqxCkMSFgNWzIHqyZRfNwQYvAzkqcl2lhiwo/HqSw2DA
TeaRolRBt2Q+6WeudNFRODmeb3fyN+nNxzs/MOV5FIGsfHcdJcujflIJ/S9vCB5d2Gksuz1Vtvgs
dEoxVZxMp2UQcjZrNrIVnF9zNBZu9AsJ72aW+enVXrlqDr6ktwQ0XebMhL76voPt3fwF2TCUH0JE
MA2H9b7U/JzsqDQxHL3TH9b6YOLwibp+ZYHzJIGr5Zq+6zaeNr3LuGwTBlu9Ym211SUWUsttByy5
SSz9Y8Hsmc7G53d7ceYW+tXlLeowGzXmUiFQKw/DZsem2ZAiryfuVkVgnWq7xGZ27QUc7SCZC/mL
Q/6cPSMJwr0+w/gH8y6MFOq3a2aG36WbaT0XDaeMTngLk+0j961/7Wajq1SjhCijYZ/zA4gQcVmw
t6YbyiIkpCnfNCu5lpi8Ol09MTF2CrjQ/Sf2lqWIGQjOvD+JXYEm1+opd3IXsHJ/s9SqeunTj1sI
OLTR7L3Z/YcnE0bNl6vikxcyMqbNV9o0laB8Lse2fymcdvOpEo1S5VxCHW7nd/XZswsXEtn76FAW
CNw2V0GxRUJ0v7JtbxoGMJXEFWy2/asnzMY633RPrB3yf/v7lsd63ek5sux0V3BkdWyyxmxkRx+1
cOcRnXIIxUGaU+yGrY5JuAmuo9XGFM5XcH5oFzrWf79zgEvLUwN1ceHUNLzSONgJjUW15fli7Ml+
KoZQ+SSimDJ3uvBeiHyOgu+1zCXCAk9zYfhH6C6YngHliwEVfd2dF2sC9fwHcpzrGcn1UiGp6cQq
i/YvxjMbRCAb+eg3hVMDQ/pD7dkYgA+NC5HY+3vW3Jh/kB/8P9Bp051qHfinsKHLhsQl7dqgeJ7m
kwO6I1BEgVRaYrj5lqFqtdukoxVW+5qw5FUFA2H1kKsp5tmCqcWpDfTD1U3p5VTRQ0/k894cwBnw
RpTNTmKjL4CgQZfCp99uUg0mJEE+13H6WCRM9kjIUAepvXHBjj+sKySpH72JB3qF5cN3R+WOd1n6
1iZAQtflDqlQc5h1G89SKfrOqpkj4m4WKn8niXdNF/smq5Rz+Ij0E9ii8rRdZAO6wbrb5MUWUBTu
YYSjy7zYBjt0YFGUrgVkHqfEcqsMAfkRajm8yZkKF1fdLDwq02lxr2F3OckPRJ4mdZkjoujueva/
00rufCc7HMsQr0l+QmJtUxapOBiggODMgy3CefzX631jFT983RvsY0lLXvol41bETsaprJxuHmvk
cA0kIQxC/73+zHoJvXb6EffX2KChd4vegqfBcU+6fLIoydAAPr9TMuU1r0mMzGruyWNIB/JtPqyx
YN9ObJASM4E+/Znt/wQz03ZZgHBSClkOC3z1FommTY6Y1QhJUYsq/fKjImcH5NpCSTKzJqCUYsmz
fcgPI3b3+KGAzs3k9bgvYTsANLV3NXRiMUhln1T0K8hMuh5wruCe2qyIb0a8zTd27knCSxKA3F/1
8ti666oVIpruan7TlgQbvOiUDzGwBDZvl+zsixD8hJt/t+r9WQEKMOae0r5kbpBmrAL/kFWUa9e8
C8oZdxItfMuLOiq3x9dj02Yyl27wAVZ4Ba6ff+Ds7/LP7pR4606i+BP8rnVxBznBo/O/Z/tu4no/
1lbLd9wUPPq3p56KQiUac4RV24OUgamb3LDIQAT6gx+OXsd15X0gpzaohRCpimWSLr8CJhTw7/zW
G1KYu8KqguJv6OfGXJIroLjyJ8rt/U3vlwidsixAucmu4N+KqFdBRjBRaM+6bjjLTblUSj5okM1I
PXxJVRFid8oRjQyUHltvp3Lu2IISAEBYWtrmD6ezr3BW93fNbpQZJxCkYzQVZc5e03g4A97f7Vk/
Hz4wEFSnUGN8bigg6vzHFDQpRu9YnRc1Z+tcU9r2NTRQ3TvWRISDdCeQhkHQ7BahYZpP/HVLn0HF
rGgsIOa+Z5fabcq9MKko+CSEKHUPZtQpAXaf62luSbmI++SJBRaz+UBzSN13Bv/3VXPtuha/4hX9
63R8VIuMjmnUt1KeQHrLbnCaryKDNqS0u5/wS+fuGkWVbxFuvgXYqjlawt0gCzJ6DSgfvvMQJ0zX
T7KvTdRxBhzIAgfOsWh632MJU6t6ZcTN0WkigeN3g5crCuIDX4Wtmf+Lx+HCMD6X01p/EJwb7w8o
frdJ0BBBQBYpxqCct3dawsJNSUFocDS2Mi57klIzlw9S34M+rv57FFVZk1UQaXUJk8iWJqmWLZwD
3Ih1+kD+4cLbtjN8qslIikhkXjJp1ybstlll5YHkJFdGBHt1vdTaHbnITdqmlokTczjZMyKOwIBE
4+lx4Wl3b5adhKDdxxXV5G+I8jrAq0/oAmm9z15V1rjt2IFChIyBu++vBA9k46raZA10alrDnB2O
ArGHEfW8cw+gm9JJ54wKY38UR3fCb8uuWcAQRYVw6lNK2Dpmx5F5xSLaZjoYnGFtze/hhfSMzNw+
dZgG+mu0pJiUwhlBsZdlR3g3McjyE2gkuzyPNZK4HN92sJ5R2ZSBlbmxWNGEnTVN+br9O2UIADhY
Sahcl7Z6LNr/hupOfKUaJWRvbkVuxCZsKVtSr1xrH/9b6YgTYPiHIt2YyDE8UrfNfX1ABEDdpOkq
wASoCAxof/RgouH2LCUBlY2jWDEsjwKxBSd9JZNJ7htBwTkIA/8p81lwkyw97Wv6sNWuaXsvQe7O
Gm6nRJNwLcieo9gyY++VINxLuADOegqiBvYUHsWVOPkElQAEZp9lqzRbdHaK1Zb2lCQ9W68Om3Uz
Vj6QtvoWmkWghTOBEQg1EZqervDwyt3OYXFJw05wn0Vih0MUbYjnRL7OJI6HzmcmYIMxBECgFOgC
9VRSdDc2gLvT3xkHf7Qoig2FXHJraWNMqfIT0x3NgVuav0gHVTRZaEwttoVI5alTgjlMmrxuhIid
I30l/Fp18yyeqv2eFC3heXmI3Fw1lP6qLdq9n3CUjOhNjmrLFEQAGY6iCXROc7A63lHk2qrNX6gy
wp4Q/CUBmfCjRUF8b8eOPj2NZ+71WPAzt71j8fHzkCzzehZicids0DVRm+Eq/j4e60kpq6PQg6wC
cxF8ubXYrIJ9ekz1TzFR9t0Z8UsRrWB2mt3xcivyzAA+/kZRDiQdpTiqHP06wCF9ac/h0hv0NgH0
S5mdw9yhvjSO/UzsKQZdGvuuGg7Q/q6mBA+/kmDh9zK27WSSGZI2nbNYf6MGNKW+h1BboiXraeWh
CSlWlrOFU3XccLWCkezMmZSswZy6f1kt+jVZZGVDb/TMzZ8SKR6URSopctQ9oa5y82ItOzwX9R2t
64kiWYPuV9PgfwiP7bOJ9GYBCgpwJ3Sh4RFKBR3VQtCEv0sEr35XZd7bgJytt0SYrDeFBxDzDLmK
G8mgj+oKh0tr79U9LwlL3pTm6Wp+yZ51MUA2+rFB+/haVAYIp/0Rak2bHDjy2zhfLuXeJGmiaxHA
IxKT8jqjGgfWbRga5QjUOnrGONYd9u9Ab2ZbuhYFLIS5mhimS6onj7KuQgYvrDB8qukmtK2AE4s8
DCsOUAJqD4vAZ2kPMpHarv1NfdgSUJienWNLve6kRML6bY/jxe4gU+MXba4aheiH1ynFYjeQZzD0
3C3q2BhPoABKCmRFtDHygxZViFmzqFTiWvoNbKh7Kxn2FNrO+OCjJ+/kCq56L0dU+7U3Uv0FYqvJ
uLG5uxIFTdnOoGcbqTKT/aB4zzkbAENROuXWnMrv16bSMhClktl8GCkgzClDfDv9xM2Rw/KZ3Qi5
v8yl7j/avatYkRAqBP0RvS6tG2gVJ5E62INJjXtRPtR1nKRWN+pxa8+vlOhYC5lowz7xjPz5LC2m
0zzbIDL/Hf6TCfGIiYXcl031Rd+tqOEx5qM0xxrVqkoQGVv1Wj9PR5KvaOhC6aSTYmp7k8iuBPC6
VRoVOTx9IEce8BgaesMi6pMC57Vk8dYGtqWNoja7FkoVT2aNZVnHhC4aZNi2AqWHWq7zPlziGVTL
qUhd+EqGJ8CFSTmaQfwNuNx9cqOHV0O0UkEig9FGPKsVS8LJJh97Xiyyq+rX393z1OEUWAyFrN52
srKsYuCmZ8itzyZSkDYuHRBWu2WKUwZo/3hvZnCfGI4GN9XVTNrXF1+IsFtxq5CJi6RRx2hMy+V9
qdEN6V2KFpcOR/mm+ztuDwZNiz5+cT6buX1SiySWQhNJxS/Pt36cIx9NUE4PZnoWRQN8E0lP6R7v
LGMs9AZJBpLcaZmlVuNBlTE1hsAV5WXm1rg7skGaBKJCdhvL+/6SrSUDPonVP9RgyFSWFs933007
e0ai1ApVRBWIyT0+UO12qOyjmGxGMkTudFDOnMQVAnnLMvlwhoximcaKCAWTcQAcNawQo8+K5AY5
rLB6HGMGGzKV3qDi8DqKThDXl6Nwlk2dl/L9nvC/Pkegt82H2ZNijbbEPuuLtbKzlNI2luwH6lkt
fkWGapX1JdO+ViuC5CtHT3ObrCkJEMa0FwKGFj9JTEbZlTA/1hB914P8PBdsNY0PbFuj5Bz05t92
0etjt6vD/oJR2qfpXwfinZTmkk1+ESkRMfHGdiR2yAi0QzE8LdptKYk6SXojhrB12cxH9AMFDnNi
Jntjcw9lrUXEH0f/55UHg+sMQ89znEyKpPQBwtKiq6inI4W2v3cc7o6FlF/xe3D9NmneDE1bYdDC
uGsnXTRO+YSKznOUWAi2PgvJECAg+huD0idJTioQPIN45eQFufiK0izIzG3kuQXKDcm5adjm1in3
nQTS5Pc5F+jWT5LVEe4F/5n7r9kOuIuQV6GrDum8zGhzaR8kkvfwGMDx5+FKJxoIHnOERENzPh/2
VLRweMGiZBE5nJW3D3lpNhPKXuOgaDxnCgIXb6UYTajQJV8SXNFEiHzJwEMNQqrdhnWRkwnIvwHV
kHgM5iPyZPOm03OdHViVETQhryZvpXkaAApHMT6tKnGZ2SQUGdzQZB7hPTiGwKz67SpCFX+M2Knm
/ZmLjBYYBY9iHRkkoKmyxodbEBS+qDiVkiStPpMt8ty7ttd1JqDHIsgPXTRsdj7MGHqIVj1+9RQr
LXgMvXcLW/vCJkBbYWJ27ACIt5hX8uSZyUQErpCndZCqNowtWuSJ34cT/TmaYLx4BIP01LvZ6eNO
hPXRFsiPZLHjfUUBCc7uvUpTtSmS+ZldWWzB2NK3pztxtXpRtsXbsf63GU0U1wneRrETHbKUKX4M
e3Y3Bjd9mTJTnsAjl0/wU6Ekkcugi6irJUaekuJIwffeUBSZK4e+K4h+RbqUnBnW7Jic3WZdb2MG
PtbYo4ko7QqhEvthtkWzSL0oq88hU3kgTekgtzavtHfI0vZSjPh/aW8xo60MQbHQrvC/LngUtGIF
msXdnjn/UdQba8t2mvZsBX41WIZduz++UE69hqWWiIAYK3B+6LdCbW000oCzlp/Z6PgF4bjfSNhM
cKnZdHKfhTzCaontUmrV9f58L2LSwr2uMabxhItyrO7oKsCIfHRNmlMQcD+sBBbIe0K5hbmfdKhC
Iz3KikC3ATiefFOHXTrrQrPdw7XZJLHEgWa3AXVEOF/CLRSqxCeOPOvjaKSXM5OgAm7+btsVSnex
ZzPTXEpN17H+vH+/s/W39UT3kpgkVK7qeT0RusAFNpV1JWouLqJeNes6ivNFDgdePDE8FlPZmalD
CwL5eJe9umA57BF0aKj7ewlVlBIJ1Qb+I68uJh4ivUsfO6O1+Wj27IF3QYY8zJR7iddDdQpL6eeF
DyruulQ6aIQ95B4MxnbL30TXimEg1XKTrmmV0pMEw9k/QfdEJCkE024SjDahhuqoshVA7MJuTF0c
r804n4i21nHzmEGmUkklQMjpOcnNC0vb01Mz/mev9lfh5BHFxFdPpzLyuisF0r8fGV3wSeVquZky
DNPgw3S7MZcdg99e95jwFOeIWleNYs5+zi3muDKx6pXBFo1aZU64hm3mJJc6tBp7dX05iT+tCZYs
4kb+2qAliRrmqWb0AkXZoMowWZ3fAkDS4g9eVFL3ygEFe+1t1rKbgJXhCC5DaTz+kWoBwcb3HWMi
7hd6E5qVPrxCaHb8t3spOj2G1GLRevLeQLsbqlcQqrlXvBkYccHYaSZBFx6j09Y/vQuCV2/aqAUb
2g5NzR3yo+K21ZVmwZHR3p8Gy6Ar92dkfL13tVZzKgVJOj7BSoVmFLnQVLQRCj3ac1MfiV3qJZrm
scO0Ht/mZvI+5Q18ShkGN8MjVZObMNF31MMlowFRNB4/ZAJEao8bCjhCJMrVagZxBAnqr3UwKJt0
YdlJcr8k7yiJ44tgZpqGnzCE81DKHdlnMFDDUqzBPUbxN7vF9GLAWwIZWj8lgQyTtH560Z1kchPd
PxmMclLAlv5nVZ5BljvIclp98zZGLFba2Y6w1Z1tHhsKsyHBXQfykCRZ/ACMnSTjrKXfehl0/6rW
0pP8b0N952ri8uimZi7y/V8uLNr5047pNHQpCaIT94B7jih1jraL/f5/KU2cVR++VievSTjmcYnH
dfaTkpj5uwCKoKjnBQKphf8bpsJlrIoWUNUcQ1DfI0K4j6vmktEfkLAZy8WLLRbumG2b3x9rJ1jk
fEjIE7nn0nfPJAcT28MJN+jiMLEinh2wiowOahCPTo0Ozx6/bs+KZ+bxKtDyza3jGfhYOVevQtr6
qMPE6j7u0iGcMikl2/dt3RCsxpuFL1XcHABdzn53bGdkbcNn4DsaIOsRgXWXHEmsS61DRQ2FPb/u
xCMUII9SjfVw3lOl7jArOTXXd6OS61O9PqoMe0fHw4PgN/IC/EqD4b13fmZr7vMKmH+nEj2vbBYB
IMqOVfscXZfvKXZmi4d8vqya6GqFo+KADBxxmuK7QPY+h29hkgbleayVAgFxSN7E73OD1fR6jyQw
v3T4epd3weM/iLs8QBT6Kng5JYEbM7kM2t4TXhFi88qLohZtoueqNIM50AF/AzM+/Y5Ywf3L50FP
qhk1hSGZEOdW+XUS6SRhA0I7utWSpqBmjkXfqyIt+EM5dZaM0tTDy0ihsYbixVubDtwmCZFblHcf
Gt6WK7cAnYGh+RVCNKYv6YQNoVBGhaQYQkwg36zN0E5NjcD07Wjgj219hYkqCk6+oSZETvHm/0Zu
0Lbi6M3M/ypfC9Qa0SnqarvYHblB+Jkk1piOqi48293nnwYbTGlbnvmRysuMB5Ba07RVPdqtgp4Y
1G/bjAQxnLVkomgTWfwwk2uKQCGcwwWOqUbCMrK2ga6zv6BT81H8IY7OX08gqD3BBs7yVtWsKR4g
4SGmvjYE+KI3I9jWvld9aGj0hn0UyPGuEANfdJlhlzLWC01y73/qfPtVUmTBCj3eELLYDDsF0m0H
SRkaHkRgsFTqYKjoy2RQ+njXtNGfRN1PMp2Wyt49n51umQUJTCqFLVwsmM/iUNMuNB2ADGQJf+EA
9tJrxV9JdnBpI9FbKA2YzrKPrPJz3/DMPEGmtGp+dJp2epOL8O28rMAdiDAV3zS0E/iiVYLN/IkP
1wX1xMhXM8TS/JO6fIJ24cv4Q6wwgPMczbx6aPmqU3hxbTgAh/2K3XO7brOXy2g+LxJikuiB9fzv
N/Gn+tR775Bk9tp0eJxXxa1gt2KBjlmIgY6KmUhQANk3k5AR5JX7ezVBFyN5W2RBETEeWL5bnYcT
NPBKmEPpXJfhgOyDCX+eYGpLza1JyvdBF0lGQjmOIzCCpRACQODz9FMPKsqBpRmITMeVd7xg1aga
iH49jIJppe4cNFsbXpdiMnBSo4ab8rbAVI8s5JcTEYYOWTbODodOtdoSQmP7Q8bDHd0vGdVklYa3
h56DeXQKHRCk1/KK1IHNexrkWIbYD1xFa2juQ2vdjN02ODEEyUUL3Jmtib4EUV5xAXJ3UXLFNUe0
QKZtFm9mIvdjgJuIZV24V/1Th9AEsIxoduy/xz3LUReg9rHzUQLPcIe6beUOC5GwPeajSbQNLSVm
Hdt0koL14hth2UWa536WNg199N/yROk4lr1tK+58pvTG4pk08ikuz60h2LIvfEZsVrWpeweTTbEx
OVScCjdfUcxSW7bWXg8b0SgGGlKlTh5wR4QvX7tAcqi2rYFFtOIHFV8V0Hs16eZmoSQ3cJF6MjzR
How8ilkVgVSGg7OF/ZsDLlLZQryH6gnnkCjHBuMwhzBd2dKzgTPzfGbOnR/cSP7CJkH53wo2MnYj
R9X0+E15SJrMmnPyH8XnmCDCAdA2/SrBzz3zj1uZ/lH9Gc+xZ2CUEDVeX6cNbFrEQ8EU4kQo9wB4
CktAHgh/Wi0esZS2PU4MWtDNHBO53zoNDpMKQqeTV9DHOAE9uaA3Uql+VEUPnD2S95Axt/rBM8fe
H4/RzHPlL5ULnDgzccHbPNef0T0KlETgMz/Hvd0nS1gsjTy7p6sMGR44RsjqfAI1KMP1stwCGliu
RYPaUG/UATZ6LXGSZi/9fF6Sxwq7vn8qfyN1E8JZFhdIwQzJ2VuOImKdd+D49/eG31MgdjsKFX/K
gc1bKgZfCW0k39/Q0+SE7q8hb8Kk8WklQeWV3//VUBCrSVrVKoT1ia1CY09rTwGAKH+G7kkpYr9R
N+60kaC2WNifD/RF5xYPl+3UpBhmghtEG1ITUS0ZNZA9T3EHb5EVFmGOM8PIhNtnaBzKtEy/KCu3
qpZ0M2ZGZMpsPG/WHIDhFavGuO/XGbv8TZa435ygXkPg9VmLHYOwXshayqc4zPftyhdZyv9iJIMU
d16Bule6NkW/F+CaPGAR8rymYRJiBiuPnPToBekks4ZLVYyZ0+982PC1VOeD0csij2CpnJ8s2qKi
Bw6SBFSWoXz9os2r4uts/2F20xYBb9nmo1UmXk3xjyrzOpsKdQs6fgCCa2gNHhGNi6oDppoj3+Ze
xFo9iYdtZlHd3Eb5KEY21GFTnPXwrVSDlq2+16wG3aPKzjd4zSwqp1nopMKkvc3pYclnRjYyS1mf
/DxS6/Mf5Km2on+bihs9l09Ixmg3kCHEcIufBRwkHtVhnKOkMYYVKDyVZO1SR9cV+IAtE/QJzxCl
3AndmRcjWkfFoD3wTHlYlS5hBaaLHJJP0oCSm4ih4/ubRozm5GBOQEVMx7Hn21OVKZX73OH1SLKa
ZgrmVhVPbhf6EPPyFwVNUKrKnD3plCrMoPBoPmlEhEyBkmRj36d59rYfzYtg66YGRXIOaqWdIDqE
Vaqg8nLvdVB9B4PkSk7jEXtd/9BT4c6KfiQPkbzCTVPCr7bUJEVR/iiW9Xo3IoxXbyr+sf96yr/a
IlRFqSdnX0o9ElDu12Ym/o8vem7yS172dbjMC6dpboFu22E3BiVb96nqOjy6hZ+3pJ4cMw5j3ftC
Pi7USgB/UeQ1XsP5GOfn2hWVbbVunABfTmSpXYBn4oS3dsuws99nyTfLDC56SPfPuApuxDAzMzcw
G6KZyUsuEY1zGliJeyjBhfG44YowSbcrc59oFeznEmmS4k4XzJVGY51Mpdsf5h/kpGEfqgxDc4CW
PRFg7Zw4JSoLMxQ3FBMhyefv58YWJg97XZeqHl/4At2fHb72b8Brgdol8ReLkdJtMx1sxPWjh5kB
zxAdy3t68EnwN/HJGZDCETFiQP5YVBMm6PvqTfvWsL7vK5kWhrNUkx4TGMGDpofko5iHh5ZXtbK/
WSuvA6p7epRpurzS2MqNV7zGsmxnbvzKEcHdMImHXmylAMIv8uJWAgMyesdIVV59Y/96K1hoDlrn
i4ih8GpZGlUMvPU2FtwXuvK7U2num3YbYFBoyL5MwQh+ulKgcIw5XzkPaALZ/4omrfqsUPvptStJ
ZQg+qjHKPAgGwMO7XfhmiChl7xd3eRnkv4MhbyUXrjw2zzapJaD4v/zVionss2rV3EhDypxW6LUR
tRqp1DLGI9IWtYzCmjafRkPfNzB3xF3XYCUGNXiNNjJySzmQxI5Pj6lmNRD3x1JYj1yN/31d2VgS
8cgdzwxBZOZOmwLn2V7TL3m48U/l9cc0doGD5EWCx5mkFU8FyYUo0+qLRBKaS511k9LD27eC4cpP
sxWiTn/tzUPegZW9CVq5DugCm1tvgaEIf1HQ1OH8cGTyZix3/0nAY0mvgcOo/KQ3bkz4P3Y2Dyx0
IPchAwOMNHTzNMjhho5O+Ra5A13EXQ9qiNaFWciwpXy067IQKXkyDaTuEqYbttnEbB92fLPTZeqZ
vaBPg4DM+1Om0MXhoS+14j3poPMgXK4xyej2i5YQV6MfowZGZn8JhTholwswEDUwp0tPd8xsewB2
zD2/G3OpzgReSeh+Gn+8vnSxXGdPPa6YlfsALOCC3ecMXYSjA2/BKzD3y89o2fPBkEWSZGRT4Bsb
SvswHvyvVOUdjaeGDiq0kFHrHwJUSnSh77Xeq6TmaJB3jDZMLFNozgJdUBFGrRCt8/EE9XyCB7pn
N0TFMMscxfW/Eqb8PDqPqt8M+CQKy9XL5jUxrz9MwRBa/o7gCEI/+lZ1xWOFdv31RWCTfv002zEq
uFgA933JRTfefgei3w5CtyND0PrxqBuwrq+Cxsffx7dDQytBd5Mzc/yiI5FKrRnb/0uncuTL0MCQ
tjUl2x6q5XWcPUxBSAHiVxwlXRU6U3F4/a+3QOweFnmOff9vTfrAJYlQrskrE/0OrjltLV9/p/zw
eEQoAtUn+y2yMANuby4dANqIIUhYfMN0G/PEHQPbtnpWrILuLTk9hRynGdl1ivsRMES4b2ChR3Vd
7VsPxVcCa0Fqx8o/Xlq19sX/k036P3E6ZgQqim3Gmk2SOiQGyCm8MhkbDpMzCsC8LpMr3hl5F1kJ
VOk5d8fAjGSlsbsp7NZ8I9dlFNLxhjHTJEW+vQVAJFOcoKJ/8o/qNNSkQ6V0OrfWCRTv37qmK/w4
7RIi5VbYzLhspOV7UeZVk7iBwH93nXiAVcHdMNkaWmk20kdKOQAjhEy8UnK1vX0VK+oP1W0lGPLO
Nn93MHdXfJbVZqq6NDt8CBMDrEv0ld6ijQwxEmURrNk6SVsBwfcx+3TTcXCXI8VJlF+vcYanr1ou
bU9F8TswX9twZ8i9XKKB+RNLi75aTQMOFmcYVcDz0CgOfOidUWNuNHAmcqyae52H/WPzzcRbq33b
elSb+XDEqyfqYDBPC3oViLQC7kezRdQ9e5u5I/NlsRowGVhVs7e2sUCG7uXPe5/3g/SVc6m9bEMu
TwfeTr43t9DQY6H2av/mAgOZSnLfhlBKWakBhkMnbfU+iLUZDLy08cDlyYvnQsviWrCX6uAj7BY6
4e+AzM4AX1Sb5RnOViKaiCQjC6EVcVOkfsErbHFE8c103d6N2QjHaXjRby0XFna2A6cdzDESthaZ
FYHRY5MU54HHdXBcc3AO2WWP910iTKWRPGimjUI6ToqrVBGTIDh7FTtogbp0L2zVolNZT/MwwU+p
8v9V+SQ+3iHgIP1r9+7pQt9bE94Ych7l8kJmOPcZ2veTqa5jIH2L1x3FNfauMSbOv+pW/58kdm27
Zzi4MqKCy2tGEyAfDI37YPMgZSK6ewnHdcjo2lFZNkzj2WWQCdsglp6y2NR6FOaXuO0ahS6ZTVUS
FAcibU8VlOK2XAke9MUpP2+SuM0OprwEsFIz4Ca/DlQYnUaa3y4vBiGBk42aFXtgc5pYB6c68ptU
8aWFMxun4xTlSZsiZMyTTGwkAtfBYxmr/iNqAvPOtsI1VhLs4ZUccREm1nLJeWSgWtJnLCmdgjBQ
TsYsNsjYtTdbnPd0lObO4/KIUzt5HSaJedrztAuW0j03koGn9IJHCA3mw1UdlMac/pXRiGwVoBux
DKSonq+o2S/V+o4W+xqaqAOKms36XD8V7ypmX7/JhLJaail3GN28LUOE3UdMx9SxzcLb/AShaEHN
TZNCvfZd6OYvlGz1r58a3KgyGgBwCx6mutZNGQSj4efo5Cmq66LC40cAFR1S4UOWgDxFPSaELs7h
+vWXcDamAuXsUN56PGOvLFFoSB8jzK1uBgOTIz4V2AAHJyHdtoVupxOYQ1zNKGjxa+cGjCp6xuot
+XsmyY4Q+o9pUoSIKsLkC5lNylsSoPeYACCDLAXKGIeGyazaDQWAm6DCJMrWmcNk+74lzcLgyXN3
WNlT9fwazbP7CRG+DGVXQqG/2evMNjy0VSak4Z730jwsRKSWGHCpqhYlKeO6fN0WP85LQclFJglX
WlQKbfdF7goEjzFbMVDazIw2/Vxgca0kk7GuQdbxFjwaqy1NuuQyUJSlRbDZrYRT6eIfY2z3zCqA
S2Nz+A9Fv73S7PjM69q/abRu+ezzN72YcFluGB+0c19yRV5+2vmxqUSIUEy/TjyXr5wBvNg1eACz
zETTBgEfa3rmbT5IHg6i55yBo4F//0r2AnQUjQi4Hw6GSdwr2M2f44BADGXmF7sgfRrblyq6ujii
rHkRjaBHu+8ydutDdHueGX3WB17GBN3h+VjfocJ8uLcNQIwopT3mA+UNmHKjCxlj0M9bNgfrb/Rd
CtHVvP17K+p/o5TvJDF5JSO991KSw9pDjCAQ320Tr52h6Mqp4ZKCTRUiR4VnHXTNfeil9LMcs5fg
BUenWWc7cOzw0NHmZLuR0mMfZ8LaKEpFop+Nt7fOQXVRkMWIuGMb8VIxi/+PudrjKZ2XJmPd4QZP
UQpvq7DfEq2a2ugQ3FrumwNW0Eku8SgCSNTCy+rUYKrhN+YoVEuk+yqP54x14OFxDiNZPfRctru+
ciGPSPXlxOVUFjMWDYM9nUOaTdFSlK4LhmadQAQnU3/ox/3JcsusY4xiD7DG508mVzzQ7/X7ri4s
jANdOx6CvAb5oTeIOnvnhQkIbts0MLq0Rq2uR2UE22i5URuFbM6Bc2n37NWOnuqsb97Goa8PYCuJ
YvH2TUOCWA0E9eQOH/oAzrXHN13tob1Fvv04aM5Ho6LcGyFmM/djoDcyI7v3Y8U9J0SsbTidY5LQ
wrJfVJd4mPshM6URRDgvhZlnsty9KQ15wSxzrzSW7s7U8fRv8FCXzZNGj1Yjf6COwzhhmMFFhpmE
05CeqHHv/jEGsjMp0oqR7tISO3VlxaoCaqKWWgiiTkBsAb+9tEQeJSu6LVZEXwA4f5aZJ7w3PEuv
G0byHB6LoDFcshVHCq3S8ozg2CkotI+ecMoQNNmEo0LOWMtAyfpVjNJaweCCZ8nkh505r/ggKGDB
Min2YcNrXHbfFKtZXTLmyuTsSn6/COSD4Ozg624M1uokUW8f542+mCeN7vofVizvC0ic9rA3h9MX
tXdv8iplnlz9vePq5QEvgqlgfu/SZbVdTtu9FX72aqMT03iBL/GQZaa8sZIxnUmGnHIxCLuRmnQA
fY1kqh+NDGtfGC+axi+uLHN42W1bNiIFAJ7J2uUX9dAJgM/BgR9q4ObourFRqziJRhlSqmsmdff1
DGBF8N9c5/g6pkeBwM/LLHsXVRjJx2AYngaI8c4JlLGsNY+D5iC1Pz25Ki1+flAIZtxfHi+7UImu
GuNKDr7QbpYvaNyYYbELVO5VX4ZvmA5yzh/yGuECntgzeJgvJLjpPXLQ/hA8yYWrTY7ZDEkWa21p
CQ3I1TP5X7/3FVL1AtCKlE09bXiuzpF2tIKlXdwE7rlg22GUvRe5m6p8RclmkCDlGfcb3zvkrFET
xp+Lc7lu7nKKM3WBuJ0BLsGeCRTVkuDNfciiRnvt0oSr+1xZ4aL47vOkqhKYOQTwXpnL30ex4u/z
ubvEWwFQwlOH5zbYI10qOixYYMc4U5hvdue3Xa2K7elf75MikzB7htKO/XKuAmK5IP91SPUsrQDz
1NJJwRVMXySMA/6a2KdCrJVXdE6LGNfKiHs3rbAxJ7eCkmvBzyOvpABKuow0guu/anI39Yo+Jcn8
8gK4RN+jHRGpOAW4VI3WHObyt+mJPqt7wYTF6N6Bk67TRKxTTR5iJRTraEDi42JFaMN81+CkwRSe
OuRaK0klSTsS0AEUnVxTaWZ07aYe7aUjn59Yofm49fye3zmF82UlNGQ/8D8nJEHEA1KEV8x4d+QF
VJr6KZIJCU2uymCHNBT45srgoZGjNJpK2aqQXV3B7clnl6xZlMl0yQGAfI0Q3ZrOkoHp5uMMfi1+
Cc54fPV6v/m6PvOhFkKn8WBp86zGvr/a8RuB8oVH6f7vPdYebRl9bHw4QGiGMp5GbmxEW7YxmH8/
OyKDpQFiORl91NyuDOzxcokJBAd+YQzpijuA/QwH/jOLNTfBh+tjGPyThgPvoUQjkzlnsN3k8ZNv
Tk+PWAba1NsysK97LcqQCDWzo8IMWYb1WYAc37f/SNjoqH1iaSBBKeF7y8KCEewtaACCWYxNT/r0
AdFvVgtwnZxfLurG3zZW12Yq6mS0+Kq/sskoUnCqkCiHR+KBghrdaP4AIQfc8BLEqp9qborFXBSM
IKIIpI5L7TkvcbD6wZImOz6g6NV0LrbOX7k5YXbEPD5ihTB9zd5ZThk3P4aAhJfyWDYFzbrThlY2
4Vs/Q0/d5nJuRj9a2aVUwCs1Njf4McajjI3bWHGUjNNSP8lROaL8Sig44yetkZS287zUya89+Wo8
akHM4UDr98KxQHJUzQnRWxml9cm1DDOOtc6EiNobexXHeoBKBM/EPBQY8rMockBDCocpLI7VgmJa
+d7b29ogPEzm8gplrJ3Y3Jx4ubpS02mLa16FSdmsA3wVTCVrx556UqNzNiunQRrijgYE5vNNYUvg
NrRcw9Y6ooSc+HXPo8zsa6MRQDYigir4H8my5O8fuzaKU/UMbA1O5jV+8dRpRdSabyvClA+qHufe
Kt1D0Xqsf/rpZKEBwTBWgP2pAyfu16VvvYf3Q0Ty8ZOS+I8SkOx2JhcA4HxAc/gbwTWCzavDyGgM
g18yP8pwwAtQbiME3BiryLNKdEsAmNXDNU/PFDUE8RvOQK/lqj+f3Ze07o7o70JbDWbhjkQ0LPP8
ewYUryRFWNJ+dMrKyzTkQi85I6xAgzIMNBqOYDevhGYIF2a6V0NQC5ZQPPU5PbPzr0KjDNMZSaKO
jALn+Kp89NQI6prR2Z5pccSz3wsfX626SnbUqm0d73rWsqY17++QmSu+8lR8iQxRAOeSvRmloz8+
AfnNGawQHxiW4X3+TDgpj4yrC3hXonjflrtzyPTnsbiRS5WbH+Ne2gR1be4+E3nYDAP0rOB123iV
vS/UtuRMI4OsmtJvoTkjG9oXAuw/wvBuseBMK/zlwDaE3upY6D5HvMsgSC5NXFQSxlq0FFrT5fX0
euJW/cPAuKHHIBj/pg6kRk/RJTdUwMXviKwEirG3P5CFP9vpZcOYr3POK6kgQUVAy3VFeUSa0LNl
ZCkvk0CTymLudZavjQXxs/qwhzgVe4E9YHpeAPKiGOuRkpPetgPvuqTVvZMS0ewQuqwPFFyz4p3o
BL5j51mlz71Zo3q02DeL5LlRdbdIyTOtZ0GkxshwW2cdKrnNKoP5YMq45IfYhLAl+q4AKpKV6DCa
m7YC/5FC3JWaL4Md2IaEVHeb85s5W4636m2OETu9TeKHrCj6uFNtOoAvGd/RAqYMUmYj9rX8bNpv
nZI9vn+D39Uoki0IfeSpsNIro5E3Mrpa+e+xb1E3YErC7m3wma8SsBTAOUC6sO6jlHtT8gNOHwgn
h7RHxLk8dG8ZHCjcsIs9HnMchurWpj1LqNQE6b5EtFlvCQ+q4za4N0Ip8pX10l+As0j//mruNNJh
+yg7QSBfH9uct3gaIH3OsVIvupp7CMam1WLpXsWvggw//RX8OaXrURulL1JIirEKn5tYqCL2xBl+
MP/pHUFV9VyM5+7KFudV7ChVkeXQc3cKzk/tHZ4W1Ro5GJFsj9/LjjsRzstRCqlnLf/AxWTgwqC0
kcqq0zJjo7DAXCyki3NCfrS/LyixNs2jVz3wy6iWmz/uz21KCOtFvS3IrSo9Fw7wEgx0/SGvUegM
qMpGRVwkft2jrmTsc+oYwVv4/4CAsDFhXtnXIrPEhybuMgm34TBH2dLqJ3CZt+NqbmcWec7YaXwg
RZ6DTZODeihYpJG2p8E5pyrZ6bCU5jOU2v+4IZkkLMj/pwEvhGLMLK/CaAdLx37OGQuj1917XJz6
vtpm4zweQNz/+afBpxIgF/AH/S2goq8Glyx+5NJOig/AH9dy5w1nCg4yqQgSQtBwtklPr56MlLuO
dRLH6q8t/RfTUAno3wzL4vOlrwecBLjNy47+8W6XsZCcWie+sxMLe+uMLvRWjL7x+WanNamQPj44
O4rFgzHy284ojoCGjDKoh0ZuHc3Uk1shbOKxeKAovIo3Ss4SwN77aygrMkG+ltZmKaoy619El47R
OvlY3W68DRRfB58vBoaNP/D5o4YK1NC0+wL+vYbdsznhik1qvjqa/cURYJT4/DFuSW5DLPFMx6ZO
LvCuDwGA89RDnOq7MGNqtVAQ9lN/DuyZG7c8j5iWbTegn0o96JKfXk0E9mpTipQPTTyRgdbJJuLx
wcSzqaFeGTHzy8slEmtLo8Swgn3wWWSfuHd6DAodeP5gnFjDHdKW1Ae3aHofIX5X0ZGloLfQVILW
WfFyR4BSZRIkg89M+1aWH0yL9rzfst+/hjuO2qljlvPovLq7P1Bzc7xtaZOTpqlcZQ3RtMQIfNR1
HoqMRNCQZrbbQNZKlUTOFRixHDBcO9WDR1CXxJp2ErGHG0RxQ7cgGkfhyxON4kHMfoMUa1EXByuR
AX73yNFH8ESHSUbLBWTlhk53Nfg7Np2p6eKhK9scFvxDn80HCMrwZ8+VU54g8/DUEm578dGvAy/W
tNcHa2H8Ql/Xewohe26OF5P6q1LK0QzqOtt6Q4bLQ1cR1cKwfpRXGaWhkK+uh6KEGfiLJeoCyWcf
fetoKng4CepO2pR4vBUuSh0JJW7oRyNFsM0Q+0sDJzDyQf2dW6GDdZOMxAxAQtDXWhvB1aO0I7QH
dLyIrcj3nioDiXO2p9/ExmPFakZGJuK7GtcToeRw8k1/bKWhMmcjvUUzA7ztmRxxoqpKiHyBzw7A
jPRSnLSH17EY5XBqDkqJhFBMKVAKRCsLohJQp3GdwQqR7CiqQiWsks2AhMXoUxA0bqBVuqVG8EGd
4Dg7auJhQXN1vvjaRiUP4OaGJ8EhT5nZtZo9Ki9HqmrSHwakGGsdHP4vzgzgU4zS/Ektmr/Jgb3U
JxWl1Iajjc960BZ2rFi7NMdoPA/uJCo6tNmHa8kHqRnDnuJx5bvwz6aQXNwUR8Z39g/xzaWWwMU/
6X90v2gDx4Au31loQAtZuVTsYGKLVvAFfKqGdwFhcr2axlHcek3eYA+895Di4lXs4N91dh6z8yxp
qV3Aesx3/n+B8Co8uVP5iHFdxn7Fvx+7zmmKFMfJtZ/aKdasacfV2hi7xMVjmpnbEe+gt8gk/sNc
wU7MhAzYIxG1qYvE1ZuL4REQJM8rEmXLKfhKqsFYv4awGi+oXlSibpN/JOOUDARpv91QuhhjCiGr
jKRWjsBtMML7imCduv7eHY6178xIBld1+RwchJGEnJ+UngZId/Jvkoyy1P1f/gsIBupuVZSx0Ha4
tdeVADdKKRgxk8rCwXoZLGc5qZq3KMiznQRpGaCSZ7aAeRuGLmYEi6iJOe5ZdIfeyCxSXmlEA+mX
/n5MrMSHhZq6A0xtGZL3ZhCkNUhlLuHT5paCQ7z+ZbBGKEebjzF9KZkumiOX0Ph9de0VAGfkkWcP
NwdAkUZcUGpdRoDDcz9HaZ3RBy+IBRA+eJP5ct8g8uDX78FO+aeihP1ugBWihgurMR1Kpb9xJ8HP
uoKOKeQfovFVXl2urZ2ltOJwC7IRai+CEi0zrAOQW1Y/dg4i3+UO8gfbN6oGFTaGF3DtH7frt7y0
S2aF+/eeaV3jK59FmhbP3iPzY0cha580j2reBD1DSp+v0fZ0/zf/OoFf+ejWRFtOf9GwTeJT07aw
VAMhlisWE6DPFzYYTCk8c8rqAhFv9mdludDnmAva+qiS/zQgfUX7/pPOB2SP0SstGRw3DOnssO/p
wFm14NF/n9WiB/9Ylb1aQPgTLWl9kF7VSxH9FaKTSvwP+Xgb4UT++xDkDhwFR8iweFELygqcSQGO
Sj5nVnzmQpyE5bt4kwPMZQj0peprIo3dEUXxpsu7QK2sEmDoujfbFLMTwRUr0TmIM6Ud0u9AmqyR
7cz9waib/fWQD07ElbUCxr0Om/gM6exumWyaKOdX180qQbOjQNYZRtSFtP5l51KPKDCYBabIH58O
LIRrKnJF764Fpq3MA91cSgGXYq7PyqgpPmwLq4MXWu2d+o+qSpooGVHxPjX8YOX+mMtstqaR1vh6
JzEHnxQyGqIWPs4FnXkHj2jp7eySrxpjS9sGVBgyYx3m7pDRtyg8W74i/JmahTKBqwgzukblglJI
tCTvKM9hm1GiodAaIHpGout3VfzyRIoTDA1KBCz9k7QeU/jroTNkKhbdLbv7NNpJzPqwuRYmSzIM
sUwx2vXtiQ96R+kWVMKrOY8CGdIVQ8av5lWNH101TLSayrEed6LQgaHc97zLqdltfLUisN+Xj1UH
F8cFk2qCUQCyl/Eknp+V7oQ553NY7n96mWFO1makEqxaxZkWQBaOhjxDoixK/UKOuyQMZmkJm0io
P6EfqrqiY39gQ7b6ZWYkNJsUvjCw1MIoLoN7w701a/kirKCA5Ra9IeKPhztpHaDsHBljGbXgVKfa
YvCbSIWP1k9OM4tMSzvljp0+nH5BaDyQk7BQrfLUNA2ZMw2znHtz5tP5UjwhzTe6jpLyMY7UiNNZ
yerxfGkcaoRCNR0kMT78ec+AVUaVaejS2KTfCJDEz2QnFYziFwzCrcugE64wpWdZdWbNx2q3sdx4
NPxE/JCAzFm51+/bF0ZM3verALV7S2vhvEQw+dKrx0nf+862BCxHnAAPgWCGc+Tl9SDySp+bYdyv
ol1gJ7Cb1m9GasVjmsD50EaHRnmpePLp0ZBFrEfp/COmZYTaKtao2HnNE1ucWEMrYJtazWF+/88n
AXs9NSp+aRnbt7WNXW1QqjdfIOX8tQuT3Hv3gtqqPqGQFEk4TiRslZe8TGYrHyQwNZ2n15T1dRAw
LhI6xsox5gr8xVn2pBGs421ZZ52ojhcPpfdbbdT13dVSk4MEGUBj6H3k69g5Ej+8L6zzZNgBMewC
DcqJhBqTONvSzPwGtC6zzA2XovUNNRtQVpOA0pAD5I2ISIoZLoKUO2/Px3yvs9aSChFwV5I0qgO0
3c7ct1zSvQPEYPSDRYcigkuZop+oDJbiS6+cTsLRgftPAlOBlqM1iDUO4ora8X2oJVJQZN4qJCuD
SZBQFavHbzjoZqNXgTPvrzt5erZHJqivfIgQFd8arCvakf93B8CfrTeI+1M1op953XwUbvh+rKBi
NChQDlOYEqRlAJrT5Z7rLa7V9h3t3fZLCNpAX5pvXLIedkPF363Sy9/sQ9DCjpqCk69X1I6tZ6kb
VXBqglBtStdf2lnhWEqugCrtcMBTjSURz9kpJqjt9eqg69+r44g6aFqcRZ7rZlHw+3Mml1FnbEUN
myIA6rGYRhc9rw54ee3oy09FwMQVZWEUwMVx44abxqPr4geRdO31AbWtvi6N+DKIVw1lyJDAxW0C
qR8E5iOboa+KY227R1KRdDoL5eoax+3t5x09fqWAGCH4/Kc3W//DRNKoLmEe6HxAs+yPKeGaMjhV
29DwBahr6/I7YkZj8jcbA2AbjMtb0Kqgy9pAWUYJHXhpx83qXVxvA+JIMl2avOcr3oIdPv12VUiU
pucp2YnaTsNHBh0W2FvUa4wT85WKYPokzBv+S5YX0z3OmNk5+U9aLxcveqTiKXpUVeKJm+PpHVig
uh2lYsh2T3wrYHabLLRFx70xXx8RRMAooh/rFROa1iXUAzcOz/75MCGlaWOYUC3YVbfYnwN0u57U
NzsNt1N9XoX3ddUUyx4tPbRkVtlTMMkgdlg7meLiIJMeaVLe8+BknuWY/203MAHWtEG8bT0CTA3d
Sn8EamrDN1uV+Bjft5y933pI88CpF2sVfU/iLyogEZF17hi5VGv41QBzJTRUppoan0vRR8rLsk3V
HnaLk2IqFXWY3t+SEpFsJWx8WoqBPJb/x+NesRInzdNRNGZxUpK2pKImVXQT4F3hmhYjQ1r2CDcI
aAJbkbCMjVG8SPGd5Y1IG6SjvOC5iTImCjmv5caYmFG6R8VByNZQPzUFxmTup9mF3Q8pHMB6cJOd
RYSnr+KxMQ5/mVB8VIhMxAi/dxQoLaOzc/Y8EDNiYhpkucxnIVVLD2mpzAZ1Qao/3TBchXaDhNMY
hdbcvgDA0nKA/Q5eOrw/E4VI3/GIjU8u3iyvKcL2S+8Gw9OsjzjS/AX3pba2TYU15PCROQxENgPN
WOuUX9Xp/9VRonTcM/t4VgA6FjnxdmF/CF2eoZSVSmX//GW1xsoiJ9zJ2AaspcbFcJemRy3HtM/9
SI8QgkFMwJ+FW5QZVR/vPS/mUXNCUqhbjWWSylM5y84VCxwAUwnpsgywYNb29tRvhcUkRfUmpsPF
sMJxo2Y/hgN5j7ChXIPdaX5u/usRpUhov2RfWSR88tO6vy6t6MgmYiG3kB3nzv6MZsIcCcD/ttgp
0jYInS+d2YugQv0ekVbErg4HlMU32+YlabN5F4slJsZ26lCRmPPGKfYTJqxIuy0yAeBdM2jeZYxc
CqNy/9xqJln0DCxoQKiEjBhxYMG73WNVjUO/akjQ10CQH1NlsZqmhPNNEie0bDPnbnnQviw0HMo/
rCs1GrkLpRuT7Gb+0ZCPp64wPXJV+3HschVqv2CQDR4QbWejP0F9E2VqtEFp0wYwgluVN9wwYQCs
VRHA4BJ9f579jItHa1gdtwlCo+zP29I0ZZFX+4+l3q4QCg00cx0Xt9yixsjY65l/lTVxvk/VhKTd
1mg5JWeXCvtCmRjqyb9OD09atyqA9tI+mJV5o0ktX8SEX5uGcXwh3QD52gbhfvNeg1pkKHjI7I61
6uvSaNFRFYsVO0aHm1Gq8feCgCGL2l2/eSwYv46M4Efgh+S1E5n4KuZnCM2fDZ6GAqGB0qj20Rwn
zd2q6XVAsod85Nfy3zLgWC43VKU4QLlxTAfvdmFAh+hGL4xjRA7Vt/viOVNUOKK+hQOSUaQ7uHyM
G0WtbO7kaQn8SYnc2ENQA5wBAkqJ8cjodJlE850JHpfC7e64ySNeHgAhqLSMXFFwwjZSSVpYYsBq
6wfF14fAJZ4wiaD9/p3tha9IAG4vRj84bh6LCXXQ4LvmCM6jmLHLg/R83OnficCjRInZKqiNRJ8x
31Dg74l8HXjV1koby4ZlpXp385nvkz4F5BnkhhPKxgvNHoFGhVt+RLCJ5SLduP2Ixn4ubtoJYutP
v75YiSe+tHbjlUqueBiyShIJyroIm4FbsHyqMUder5mcAm0ygZReInulykFa+L/0hyvJ/D+C0T2V
JibyzAAHSRTo8K5q7avz1BMqpO0qm3CbMIBGoFssWcr9lHcfsiXviNe3MtuzgBh2cNny1E8uJfHU
HQ0n78VW6A3CHB3DBnAYaQuHkEFwyIfGmYLZIXsn6JYht4TogJzGC84OmaYOnrzY7Ex18o9+RH7K
5YLL+esGdrDZXdbmMipz4Nw8oBtSVdbERoW/3qBf37talAI2i2Luf8dR6aIlMPeWErT5pe11dpNS
FdJgji3pQlN9TDKH8aBqxJQ/V/KRYrL6WzIKWDh2ys4dn9vv0tBwdhi39xDyo6w1w1DxOeR9w9Br
GjpG4fqCTY3cYoTlcuum1dNXtps1WmxCYkhSkDGJijPvKJI37+WEj6fblN04hvl48YUbpr3KowyV
wleYziTXBiTZX0Gh24KJfw/YV6YQlSqv2sKZUpgkHbhPmOW1Dc2khqF6H4Is9YmqvJmls54crF9k
8TgO2yXW5u1XtEO52Qm4xipf89LSBhhgmDDke2Gcddc0/p1m1x+uSdoyNw5q2iIBLYsf7zATH5QH
CqZlv/7znJHY0tEytDhYlKxYLly+9MRd4q7OYVrMdF3wUhhUdWOSFR5goVHG2Wgbl/OgIQy2eD2s
3KUWF4mHHroKLZdLMSIPpB7sX/JhkS86x+6mkNvdkYrbZmzb3xpdu1oMG3dji4ejA9iJpFOko2DS
SqCNeL1ho65MVhrD+rrz0YRTiuoe7bcnakHTrMTP7gQdSGJGY6d20wtsrfLi/kjSv4NjEJci6p/l
i46/ykIIazULDCnNy6P7UjVjxscMnq+dJOEGCKNA/q2LetwztEbBD1aCBDaBPmjM99TL9glbj6BT
3dyvxX8BTb4sJWJubVmFB86ceM88l1UtG1r7mjqeAELumhVqJXUCZtuclaFDk1LxX9oiYqRCxTNc
ohXAR3uCQMp0J3GtNSN72AZSMwhpos+sWosiuO04BRj4ucxW+53wmKTPQt57b1/j0an7Cuv4cIjB
vCWriyAlO/4WK/XUGYflrWscJX5IYBkoi0pkL8eZ4ZwPmfZavg+j9cQKS94JjcR0joSsSVv8AI9l
Vr3T/0so0EtRBaPcA5uWjpsWnW6wfFB5VkiFCi9DXSJtK8HNHpOBfvu084XsgZIF3IU/aH28OFWD
LakBmCVmsYLvddQE3K0JtNoaglpxKF09+M01Nrb+XzVVIRGZBW8bbttsJgLqdBIRtSAEnt0BE27M
B3Xhj63OMTGu50MbHa5UarPnp7M1YMyjjwmu1pHzJoDrrwAmaf8z5JO6qF5SnXHrHtUA9n/IHj+P
HXu2YYFGTDZvg/rlYnzQbHi8GK7BP4SLGD3RVvsRaUaCpSEFYnGaw1fitTBvhibIUJbPjplwwOUt
UqaaSk0D+B/VDVcGSvVplK23oRlC/JE6Pm8gPGnru3pejyBb5oGRvatQCPpLp2ADoT2G4+LwOMC6
Rzr0sLPvgz/dCu/PQ2p+qfBhmTIU8FmJoErII0R3plFd82X8zQWzDlSpIEx2bMyDT6QZQNU9iir2
FcTBiodTydsfQhBxEqvT5EkSTHWWTSLk872g6tcweqNniQXiGBagguwL8Gzn77FmaYok2JraXt1W
0F8vpwrdQJx59FmEMtVNaYgLyB6Iv0iANayFA4WU9UQXGLb2Qda/e1kiaTXrE0SgWebnZYpuzLnn
OsFikQ3TAu1UWFGUzcdOkp7OR2Yp6DMoERdyOEHeYhReGqa/cuoZ/cN4HdYsnJMJAJygtnon2948
Z7AXfI2302AKoukJaYpnezyMxiqwkelVZ+dpiqCYHYNoYyNvlBIav4JCWWsd9lZl5w7tCrjWNKqc
7V4iOKvRirTTn414adqdbe34y0z4pNcoiUguissv/zGQsWi8M9ImkNUfRHUkPGkPxiMjnbMopyfs
BFAFV51G1J6VuBGgxkDggDjUcAJe0pRsB9owG4OT4hXCdcvV0Lohcho70BkaFA4VVG4sLrq6j19T
AZSMf4X60FDvDsLZy9f0Fn4hB4PTwy+sD61T0MPZyAPStJp4LmFmmK/lsDRllHY+oUtKpEbHn16N
vpfu4hWgTbC/75U7IZBj6A1XB86VuxXeyDeFP+cMk01y/fNDTelSuhWsYwQVgO9tZk3JpRhn/Xjg
mmqHsyzQ/QlhYr8qJXOv+Ai21wZIIjF+MslGipdEH8jQmm84rxwF0W31+0lLMNOSKTyyHWnJ4yB6
QHw1KvJwL7ie1DtiE98PgtHY+sb/lWjz5pVcUlZOiB+A5+IyuSdhwknwsG+R3CWacbHWxBhRpode
sOd69tvkyrxBcR4DoSW7/PkUXffWdlqgdYcgfDjdqCtM92xwT/62IaBsY3puTUEB+kDjkbWaAcYK
DhTYDJaKStt9yr6flLZOW42jUDwCJ1pZI5CZV2UtpVUNog3Qs8FIN1pnDvOXBNMlYF0V0jzhr3lI
eO734eOAZv5hjzMoj7x+K7e1TxUHQ8eO7K+G850LjFwdVHRi/ITgQ7Le5Uf8GoRk2uXGprdTC7Z+
Wjnf/UPpA8islmdwJBvl6aLsrj8oEbdvlFU8tVGy7yK+1xImb4n+VWr/ugYtXpxVnlFGn+oSEG3x
+Snvjz6vFFejm7EJtHGUzJA4gyfNzXOrA88giJn+mchp0wg3YwP+W3nviDH+JbKL/tQB1khAeEuW
btfY1KbxCK2tHi9gZsPD5TnMWvrCl9Hrp7RniPkPQsMDZB8Lw96PL/qSRlaQsCXfa/h2DAE2D0+S
Hfqp6Vso7pmF+VavKKFkQ/elSuIfqBFXr+//68tZuZuCMXWO30v6k9fJbeG8UkZV332QGiMRtv94
h0XrO/tyNcG9UNJlwAWgmW8YruyThKhfQd7bGbEOEJX/zIkCwzXnqQ3vpyKwHf1pgtblZ1sT6CSA
sLMxQAR7znjkZGYXJcGlCAs6tx0Xskcwc9EKLS7eNIYQgzn7+/rGpONgyEem4pJkhz7veHSv8w69
r0c+RLFqCWJWvxdw2cjnAgFlRKgjlnkBA48GtkCuKlW6w+ir/F8RLz90BR+1euGIfCgRPDKFLnN1
XHIPC6Z8Os3rymHeKgRhz+gspQPn2aiDPxKubNan0X2OUwLLlc80lmywkzhuDc+Hl3vGiADvI3Ca
fI8iIVAHS1r53En/C0MmdloQyfTevt6vVpOardSvnmpNBpkyE4xJ3B0I/aKAt/TWy/N91+gUscQw
k4yOzY1NU7PUBtf4LZUHEa3RgE7hvXYkAUKUiyLlXM3cqTqh6/IY6xxYK0nOFOMGuOW4eZuaqsuH
q4ruDPJW5QVed9nBrajc9sn7wHBUEeurWDGIeU1euos0KbTCvVT7Km4t8tLpKCkIQhWJiFVicz7t
Rh84PnwZ61Y0JM3934DCR+SW7XQyFZHOyjlhDALg218oc9l24OHpdHIXsC5n/p38V8WmxP2G8sWf
irhLtVoAn3rWbrZT4E1oAdbEOLsm0oppcnF8HVVBt5XsPi0PdZAspRb/kQ+8gqau+Ltoi25KvO6m
FpfEN/P4bxEB3IAtPPxTaygzyVkX4V+9fpPQDBUOXlr3h9GMTtajFNvcJMPx/jURV47VHJiUcpGj
mxuZ05N7BCFo79iGPudb1dfglEJ7eL9Hkf9jq8uCjxDVPTthq9bxPIb7TpT+2UZIO7XYDBMgk7tG
r4e4jP3wModjy7qEhgo2rTc3tREtOsxABf5GkwrcEzyMlIfeAM3u6zme2KMBn/wSBfPYT7hLAPwK
m+NMDAvyMt33KXAZ3Jid9N0CL/ONu1TrpUVjlvFie0qVI3DDuUs1QJQUwTisfaMZpBlykrJVq+yU
0VqPVxR1wIgzTqdGIOBL6FzmyTbIyIzAlSafB5jIIvPmq30kamRIrvjxtqrL+HeHNAx9qQm3gEQC
8lZv04zdsKNcZsB+eFdoKYOEeP0OANMW7oUr6TjAGdotvlhJeYEkghIaG9q57oVmQnaXpxiFn2je
4rqkv8L/Y64dCz8MuK1lWAEOmHIdbmxqtpBMlbw1v9Y3LEIWfWqMaXuBgQqKeLqVC7iiJeXB43LT
BCu53ogBbXuT2yq4A+Xdm1RMNbxMQWb4GpQNTmQqqneGeT6KzHCQ3/ziQEdPFgFhrg3RIW7XaMiD
2nKmc0cuxRPr/7w0O3qYJp0w6eMD+bGNsK1+X4OJ78kmuSmFhwACbl1ofcHIkU82iJDKIYtLWvCB
U8SgLdeVEN63akbrZEmwMDGu/KIYyT0lUzNPOI8yBiPeO8/3LGn6p3MYIlPTAZckGc3ANmJ7sgpN
g4ewgFVTF2nVx17umvTqVc2yEinQj9kfCc1qT1nsbEZ9Ph0mx9COZIU/5ESgANCg8ki5TLn4i/Hc
XUUi3VvDe9NV9e7fOdVmCv3i9EGLWiXeNn7JzjJzNaTP9+BW3eTigxi1IvDfi5LukalmVo38YqRy
E8M06tlU3cQQUmsA89cuM/9LtvGbQQf9z3RqDw+Ewo8jl81mI1c5YAZiJTn99V4fHnrTG2wuRONj
1L3fwnzKL81jHwgFeBz2eu+7e4A8pOV3gcS6kirTNywHuNcEgCcWLjoGp8TEVbkLwPn/UX3LUUb8
wQgMgAT7+uxZqTKEDY6r02VWqpSP5vsgHVnxrL6x65e1XYB/OC+LJmTP16IBNHCif54Jn4QDi8MG
/Bzpamzfa0rqP5WNg0Y2AE1Eqo3qIpj3F1OcB/WI6+9qivtRrn9Rdh4zZs3EaTaiJx0K7y2Jzzq4
zdtqtNTJJa4CcB+oR74c6RmC2nDtPCpdxh3kssXfSwMY/MqQ5K1deyPy8MSUnDg5ebrnoEqPjc/H
F6rYogfDnCaWyzPgUbGchUkwg+mqdK2GUzuIfiBFy9oIGKQ7l7ITQ+mHpqPxnBN05/P28eC0F0jw
JZTXP7pON78CTfu3Di/uzTrCrF01UtZw2ccDBZNmKGsptiWY8Y1DbiF3rZnZapPgBditHQmoFEn5
UUhizGO+GRz0+6RKMIsMc8rt9iUu5R4SIdOS3E0Qtc/UrQxZPfA+5OjoXQyXw+ukUgEQD0jLwXQ+
p5sVNOAJU/d+4wN1c6GynkBEuboWXebWNcX/AGHV2ZxTokfjAGnrB+iWRHGAdrRqtbMdDCx/Fnmk
Ngkm34JA0XSNxmXzWSpCIyumDcw4xmRAy3iWDeaortdhizvpSrnmqv/Tn03qyIf2sZHlZhWRe+xo
VObvE3RNXGOrPnk9LggXbDceZ7IAlGENeSn9GKkJOGZRYZkQ8lVzSEj1aC6mWcM5Uka56jjF6DlJ
fnDQjmNS3HMrTsJinSXSUYmbsdmMIO1oLn58wWt8QkdQVGAk/hXOSe7iABHmdcGKFSVO8fU7q68A
tCLlul7j8xxoY+CVtDE4ourgcPkkA8WA7ZOUZFbLtjozGuksKX23LDETqGAKXD0klJJOsfZRr++D
0kvXcxCqDOT/geL4JSCck77RF9DFRRfa1UWnBB7BInTaORbY0fpuX9hoBBv66u8Jvw6ynX5vzG5w
muJKotOyCYGFL4oY0oS7Y0EmpI3P04fC5WPmxX03YCB+qa50BfYT4zVXinujCiiJsVGyiUkPWWe0
BLgN3dCauiDIMzGSckoHyXfhnv9vhdCZNJvUK00Cj4liEldeVps9dkJWFvvIz2UQ4MCzZ8uCUoaX
63QTdOcfz4GzR2ItBbnh4lu/7EbDhbC1wUq5/RicPv/cwr+rnZRIwwMm9M0q4Qx+rglvHdahb7o6
swyBp2Ku+fWwEhkwzLmS3JlG+2HTcfBq24us+2tyAV8aQB8XPD5T62pCzKNz4Ie6O5uzDq5m/4Y1
eNQEoOWCh3D3+Fk4I5Z9D15PgXp+zObl9ekkIces2DgXadmpY4iNfMd6ysMAQg6PgLLeNAPMVKG/
944iAmEBKA6lo8FZAmM+rOUnDlS8CggP4rGJSY53BFrG3WQKyV1rLoS27Zu/L7ogrSKTLLePGjZm
5miySckUu4XMA4IWY3pWlKA9uapdHOXKIbdNUdWSmzbv2bOTrKGI+nRaFNp77n9tKBfBA21+ocCG
iIYNIecDjnCKFSEQ0h2sLdBKorFpvNUvChDQ9ZimOMHTzFRD/Zde52c5HNTc8ZHbApRsrsOghvpg
fc/jjVCE2f6AhL6nFHn8u/oSgAxv3RNBYvpeKubPbb8tdugIJUmH6uhkLkSHc1Zkzttc2vK/xy89
LFOg6RPLPZ2HFIrNbim38IyML08TKCkgSX3qr7OhkzjgpClK2WetIHyQ74a2cD/jSMNxIHJAvEOH
8EjChGoGCzRYtBnMp2YUj3H/yLWQ/Ee9EuPfCE6FlZqyIXSrp2KAeMxN0q4Bww6D1WMaOnx2QtVJ
3LUPgxlEb76VY8t79/d94BZOhjYJjTmLdhlnhjiD+b/CPKWr6xJVR9M32CCuFPG0BL1Sl14PGg/i
x7DxRn0TL/F5IWRMtOVqx2amItpC8aJNsJHqyT0X/KNk6VurC5A2Og2pTNcofgCJx7mlkCF1CvFC
j/bEfqQIQtdWgplrCsCTemfcIqp2Hlhbph9JgD0MP9iZkxXyRLTNFJ0DqYV/2J/jTb1lcK5ylf/y
l/1opvDI7KuSTiWKN//d6NiGs0LYx2Xvt+HrXHqt/DX4jyuFqwV4TTdkEj0Pf5Kjpm+zhT5JJuqi
qYMY+C4W66/BmQo+p/4elly4e7UPh57S2cPi4gcCKp92rgVlhs1090fNIfav4ATjQElee5GhhUz3
Zb7rh1k5O2D+qlBh8dwNrvVzanw5PJ85puv7vzhjGglfPqnhEadXsK5y2JMOeLZsZYgwt7NYXIlW
ivFzifIlqLRLSfsxrrtjYtXlTpYPI1tLSyvsC3T3MnZ2F53xIhIGSnKDmWB+bg0vQACKQ19gHzw5
NptaKZA+L9THAw1cAQW/wDqnyy89EjUMufMLRuomFkf/DNNHDh6ufzjd7PJr0XRhJa3UjqpTvFWG
cOVmU5ujP8rM1GD1TSIyGfWR5KT87Z+He58r+ogHMA+5obMK6up1L70YPOoDHZTVcJdPEAbVlBEv
zMgDUImyXQjF8M2xtwCPmKO61g8iY/qjYxLF18x28OIIu/omaAk5aSCpYXBFqG8xjGQ+On3GNKo0
IZMQrhBp3mMes736TA2L7OuykdKn83g0oDzLKTCmxi5J/o+2N+XVfTDcKhK2SHDqTvHbCFJVWCTH
kA3BRn/rnu/YHnfkomqbXpIwQNEBb6aGthicZARFyYsjxBG3Dtr46x2N0rFiuHaW+RxBronVmXdr
llWOQDEj55slfmBJqauaDV+SDuuJ6Xd2SoGFvN4u7t2bToWjRokKvqz/zEw7b29dn/dmJOu0xMcZ
6+BQgDYqY3Jyozw611q5CLjqdnGVDpjZTcuQQLwX+nlT5phaBoje9T5RRZUHlq60QGJH/8k1lpYs
vziieRfASv7Dar8gBtcwUyqGGJ+LpSJonnJAsGfFrdi03KcEX0YiQNXUAMwCt/wTIS6ptv7vN6R+
m4nc99KxZp0O6SXb7wvjuGoGaWdYywie65UqihC8pGOkhzeR0rJ3cSfcj/4AI2iDXWqFxK6GML0Q
+vvuuFTiqXK2nMK7keORTgYSt3V1tbZ6XwmwawfFh6TOAaZuu6/eRsL/feKKv+ELLYOilfX4KhNW
77q6Uz7lRztNTzURQJMKxAS/ooBZFBS6dBgElzSTDDvVW8TQnYDfdoQyJPoeK+gjmb7FHgWMSPOL
OaFQX0OIEdxua+kTiAvA6lc1lN6o7mAXffFfUx8a2EXS+lQpgF0YqWMPhv4U8abW2HtTBg/0WPzB
N0ebtRU71jvIW7pATqcnG0K41fVtgYQFNkQmNUskAq7EZyM7XDyCyItUjXKDsYDUbG5odRF/iNY5
00d27KGRqYZKfO8Ts163dP5SeMP10fTEwtJ5jIWiUf3EylekSF4BDzNgCO2r2AzZ1FbWwaSaCxg1
ieASjJ9/Ce7wZMhXfYSi8vy53XPTKT6ngOoaQiZ2SK6meQ6dnR3gsI1av24+J/rHJ/Mxye5IjxUF
LerEEjps1Zkjg33BhcPECD0pIDOiRXRioqyWIyOLbXr1k8tgeSKBkfxj8FlBhtA5n41+6/Ot1e5C
uh7c51rMfZh2LbhKxgUFsHzdxpxqc7ZJdUIIxP+20rsf0ziBiS3O3rrpmb7wvbXNTqOz8PVUQB9S
1SGV2s5QHsB7nJSiKeTNUKFvZqfxXXr2bQv7Fx2ECg0SY3rENXB+Pzxs1muoC1ucTlE+/i498PzO
bxoiAXRIW+lB2r2brPbJOqpPoQ/u0F1PA+n4hzf19P0+6apacxUAsds5Y31fYPpKhHXW8vQXKZq2
vnMVb9hz5qYV+EirMmc/UJlGhsOyuj3qoqxvTqfs+aWEyI9/D5OTAeyA0M+9zIP9xW+N/+wdGCJ4
+i1s1HtrmNxApRXRZdjQ0UJmtvaj3dfLIEt3nOJw6u7W+kbWvL6qhmjvZhFwk+sJ+w3U42N1zWyL
XcqNJpHbJwmgCgTb9syF0wrUVp/+7hSvABVuXbPLIKcMkFu3+cnfUaEsdHNc+DxRq+1asvw9PCOo
N2cu9axTFqlqj6Frf1M6BYY9A/Q2H3K5lxEdBOvwmROSMJZFBYXyGyzc+gBXjhy14RWzAdSd3Yxk
QesFE38i77K98UbswgytFE7rKD7YUBapIUyLMTUHBUHHxDYdQX7pwM72B8+GbftyX5xryhCp5MbY
Sir876LQmEF05ZppsuDgppQOnz3oKIzF8mctrKQblM51lHHDq2r2lhsr9szYl4b8DQ3XOs+sFw3X
ilndefNGPnMBqwbYEjfmfjlDw4UfjW5KL9sfrPjkDfv3IxNWu1L2JAYFSDB6J7KSY13g1QYN2XML
ukNiRQF6qTMn9YL5l+5oMm0sWiOlJ8EDYDUm/oH8Iv8l4VGE7iJjXpbm0l++fPQ8SCWI/z/h7Jfr
xumbbSUAwl4yie9v5mbmb2pe9aJDPT0xLK9laQk0L9+iQWQNn8rUUk3jlkKMUFI+b69zivL8o/ar
vB/kRK4B0jkO7xW6P5bt+zWRhOwnQhnI1agWeBKZjsgrjt+xzfUo98okSvakKuT08uG3jeTNYWtT
huiDu3QERT+KGWeS+MrCiAVd7HIpzUhUNTD7uaGtolIGV8H/wbSPZ1cY8v4IWDH0nutXB26DNnV9
McNSfgQnWph5bj0J66CSv0ycorn3CpCsSa6ffEIBOWwt6ke/lekhP53xSECs0mVn5OgEmDD2BVXC
CkNkUR9GZidocdz+LkbO2054ZQu2n5b12B90tvIGe5i75Cf4kpUUoH/Y7JiCUNs7il/GpLm0tS/T
QLvt8sEQ3xC4gkSH3qoLVQ9AtEHXRVmVoQiMMf0mZ0/3KzryhyYsNG7p1pU0NMCpnnGCNmUplOM7
yvg2Q98lj+IDD6J1HXiekLVaq12vij29+qo3XzdChkUvFVdugmsqVpm8T5HuN+6TCCo8jAsGhzm0
bN9umrZC5csd6KschpP1wgBp9syTnDlyWjPEVGkzOElxfWtyglxw/WvSMrZIm/JU4FLh7swCybOw
PxRcFMGBobnuHXEz2paPjmDEKO5xgmNS0oU7uvKOWwfDPEYKFBcMeBg724gDtOL759xACQ74AHdP
sQovqnKr//XHLcZLgMh4MP+Tqex1ygTa5gSJ0QOXeZ4w0r1YNn7HFO7ZjDTb1dNFooSuA5VfNPIZ
gHXNJalEvQoxePU/mqCgWnwKWTmW00hDRVvrSt5C2hOhoIzVRlORlQkV4+cMlheHhzQpQveErO7w
PdwawKNW/YiWjUUI7StqsdZ37c6GYdF2IRaSyJlBDj2NCZDwEOJKmtYyVmr/iyUBEMRbecv5Sxjn
QxG3ubUaNQFA6RhrCh82QOOpsoBQXSQjFTOVAhNUiFMBzBs6326Wh7ruQOBMOqz3lx1loEdXPHPH
fjD0T52pu5dm4OJKV0SBhWngLmkAG6LOPYPeD+QJVrZNuTmV2npJt87FPkQjxfUeezV+WpW6IjJL
O02csb9wDKsXkRWUiuKwyPSXkVAHeZj5m4VWJ8ok06/vKRFKII0Uf0jLVXPc7Vqjwt/wcsAkQ3bm
6iJLj3I3MieTfDW0XwcSHQPblSn6484pvGBwyxfHp116S7RPGKkPXV+ezeWxO5Y4t1nsFm05giMv
NsgviY6/YULpu7wTy2NmbrrKZQfIwWRJ2G86eHGPZIqEcJCHWsDQX2/LBPXFtWwv3vP3pCV69Zf/
LyRmO+fVBgSiUzRogItwzd70JOMJNkJK63H3n+DFWFwzdZfwUdEh+EeJPjM4O1lOeeMtiZG/i774
aA3VFKGgkTQ6jmTtdOddVUN3oZBOLBF138rIiwCNQ+eZDC+/ZIPr1o91t/ZeEPoyV3ijTk20hXA/
664otUTzq8GcR0hNgvhTC8xOtOldZddX7SeCFJYQJdcNiuYB+cqIBPLJ4LfaF0NVd5AVO0RQY+Cd
+c0g1avJr8ZONttGYERUf1im1yKQ4huSoEnowP8a8/yvHDAR+EA76K/Kc5Cu3bFDrDeI8xm13+N8
Cwdq3DSsa7NK6hEXHzoOF1IFNU+iHQQE8HbMhkR0bWJ4L3ejeiBR7mLT9CoBBi1n180UXAIxG5bX
2alyPBjww69MjBeXlYalaeUr8KEg4nKUeul5rmShHlG4kGcjIc9nfAiSAljoSxuX3OAtlgpA2D7j
q54CHi9+uKeIXzyOHoBZxUtYzQuelS2jb1x3KuCbC+FbKrBHXhAEKQnSEDx+DM0FzX77hokCPBA6
7AthR5A9oQGE+NaXHQpVCbWVk3Z4VWreIuR6hkTRQJM+Ja5yYn6g7SDFHcm4BNAer+25yTK3A7J5
3GJSvKTOQQ3+RQ4x8pi2i4sDswJRabzA9PnTpaVD/PDU1FEz2lVXJgkUFptuyedjjcv7dTzdk2+s
rhHylttgk03DK+Fa+zFvyLNJZwepzmvDONYmp3jLFF+HWkPINP4pC6IM4L32EXTaR9kxuRcm8DyP
cJ4jvg4VsXIsMuQYuAlA5to6duUodrCzuGXhDKsWY3kThCWh20qByhxKGnAhCMqSjlyEvSLXGeF5
IaiCrhkCIF2E4026gwSYOIXLm8RieDp0K+oGgce4018pYKeDSmF8PRRxickyH2ZKibcPhgUcyIb6
dohThD7Idv0qvmy3YfQ9xmd1wXX5QmoyRPMmYParH4u445WFBJtzJvmx7GHeLxzXMFjG8JWy/TdB
/sIRbGKS9ZRhQMNmZbJZn0G3ty9CJ+SaXr2Psd/RTTP7CMjyXI8UjkxVKuK8/vQm1fhy3WnpJ8mF
ka4jX06dk0awwqjHrZ76Z790aWeq4UJ9szaEZ4tk15P0ZYgSFedsr5dxHS2/wZXoajSoHkMV69ZW
7sB5w9q48BjhXEx2YcNgvqrmOTWndXRFuounrj3JeovTYVNDwZ36CN8sFZNQtVoNOJH+qxP0iU2A
o9qMzE9i+wUnBqVVbNJBokXxCv+2/rNt+l3N6AsMZo0MN7H8SMl71CvomoB3XgBGXw+IshaPrvq0
ftfjRpsBG689NoEFXjnWmMuYJqc9o+70VszXJcZIjf3x9/voJSsEeaYjCfDsfMl/Rdq8iuqVov9P
yd21euG5n17V9ECGd4y5IL/PUnZvmyk15S5K7qGnSmtNs5MqTQxQyzvH6zhtgPuIpeCIF0sneVP8
XQtF8ZpgomZflJy9RMQnE04HlNK04MOetkFGoDP4/FGhRJLHZy0LhYMa9xp6EA62PWDchovkXpXx
X4K4R6EGOd7Ze5ci6RNaqBHONHLEeJJhuILmbYWbMZm0PG1VEyDYh4SU5KXV08iJsZLKoAy/tDEC
14EVE+VMstNa7d0jHah37ZnjeEFP04Qh8NIYg9XaL89u7KHDR6IxiSKVYKdy2AUdPhOxGCNgXEn6
2jEJdcvJTs/TST6WmLRrb+Hb/jb/7FO2UP7hn//65az2npCcrDX2rwY816GHYst2ReTebIXyQito
XRJgnFbVp2qSWkNrcX1zen1QLInedWgcbQkkzd7a4urw3xDasDFXKdOK7XR1Kbmi+Hy8Hg3fNZvV
+yqVsSTCQj3sKRxYl90BTIq5+ZJGBO0By932SoZIxxyO7uSVoa+0TnCkEBr/U6hxtETSZCwNd4GA
Z2KEyjMT7ME8yQfzJd7ghv5kv7yCkN9G+xbIBzxK5YWwGSUAtSQEUqc17b6d8yfA5sqrN6PuesoQ
1PW8FMq5pEKr+V9RLV3E6Q1bJtaZvH6TJI/33Ntkgd4BmMy63KTSS4IBmvkWNUX2p1OlWjZkqL4i
scO96iEMA7lIeJTg5vB3IAcPqCcs/GrKelaugjUc3h5leyyA/YThaFNpHwYuJqhyN1AkO3JEbaQ9
0A4WJdm/yz1vxC5aY8VC5YqD1GIa/O/SB4Hm49rhNFfU95RLs+JyONgrl1+SvU5r3lzEkSXBYa9s
D+g4/Pb1yUYnMNoaEUrN9vYyKpvoPml64NdhLKmNwWHdw5GpPZ/siH2pgGkuwjyL4lhKubbXJbKj
UilonqbkPFsayjeXWrMZuPN8JvWVhf2qJloFpaccKk8xVzdhEf8Zs/Q4D3McOhAdcsoc7ZH/4pja
Nl4qOV6C37qm6NBAt63QP358r8ucL4+klqIRCZGsx1TtuIT0FT6AfPNFd6A/TpcMRdWYrr9Pvo6C
6dvUYXzmDYYPhDvTl0oOyXW9ET24cIStproAQ5CyiZZyMPuqTl8pnfKXo9jA2sRedh2LKKDLUibp
WBLtaJcu3HYCEM34TUAyCvVowCdxHRYFgFHoEsPRf+psl05HdQ2XONfWwYnyH0eOH4N4TY38Yum0
tAz14E6BOoNR0Pq1Z2Ngm1lO1nmTTsrIIXPLPdiYMHLdLK8NrXrDJlu+UHgJNRLWzKI4k78FTqV8
Q1VzJXM7Awe/xSUyALD5AlDRMr6InRcoz7fzgPXnWuRYYb6qPiBHmitkBRPIyHyeQrlfa9AD1e3N
vxluN/pCi4UNsaIYT3D8cnBB9yS5gL6aSKT5tz/4EWk5Nfa0duHNJwt/XPU8fZkPKeE/ANupeVDp
T6iOoqfvjlwc3jn3TS3WOzNVhlniiAZqvg41CM5xIh1TkjkbftUsuogACiS+oGx/c1EtDFs2jN26
eJiw6ung3fwIaItVhokiCl2B+EhPs5iJcgoQt08wk7ANXka+Udz8VsknsGaiDjX1IFlHmjAB7NTv
3OhrQivUg7v3mssX5utAm5t1bpiMz492mu7zX7syUDghGZW+4M/oVcqLnlnbvL6fgm2O7juo1+vd
U9CjauqVZoQ6BCXzlO4Mn+JuUvccn4i4I4RauDnoa3AA5FoK7VCQcBi8Iv9QyW9s/EG+tPVkcdAS
WDBjd2mtBsk2no16cDdt7Z2ChVQiVloqbQem/5HeRT5SdB2JQQYYLz17dfnbVS1cwNo5Tn/3Rw95
6iF8309Woh4ai2xqKDlsdSiWwjYNDBNUrKB0ppVJG7xjoEJOmsEmiZhiHBhDuIVSzbB5tAsBHCy+
cYA/D0GH5g0Tke0qiTolgojReL+4nloRvwlFRsCXe2QxakeP3BURwrX7mR0KIp9j2fs7SDfmKxZN
E+Gx5fMELfMdV5iQJW9H6jGHPQn0XzY63JqhE+V8rbk6IxosprrFjIhnDVdqrj11kI8At3cg43g2
vnSGiIQjO1g8iqT7sdUuVX6KVYaBNmS+vF97+k18x32SHMs3c/O1WQ48E5t2eUwTxwuUKBBWAe9o
e+tMT7ViWyu7ykPOmMVu3mlQBK5B03J4Fy4Pz+IPWgrrY7e4HUEcHuOtOO6VcoecpsMHWOAJGw3J
fz4JEY4LUfgYmWIS+9eNzHtMi9g/zCSJqEVmhcrHJyED0BsCQE28kXUlCkLsf6sY3owfe5WNIZWM
kWhaPamPUwGTjliqAihgk9m82t2d/E1uv3ukn7RRcTpfSfutRMenE0y4tQb8ydg4GhP3wlekqA/X
miRQYWQdQzLMpoajPTmPT5jxW2f2K9aFFKRm8mBXwjCGddwz0uC4/azqcpHdcs+WLH7/YTwF4/CB
o8Px9O9/kw5bG20/sOv21qc3xnjQaciVGtVZRUKwpwcshe6a2qLB9Mxw7KpkSDyLpE9IFJ4F30kO
Bcl3CVvibi9jMeGsqVA7PNlTEgh3MY22ObT2jSGyTKv0RMA+MzpS8XH9eWR0UCH3vrX6s+XtILJj
cchkFvj77SRW7ky0F6WH19i3zaAwpXK5V6aqcCiT0ehgoAu/O0kduwMTmh7Rm1K1zO75jdKUj1eR
bF+IdMtUZjP6sx1VG8lhaOUKq5RD4Uc64K1cFM2vKy3n2gyVHiWdSacU+BjVFrh9t0cmao9nwXhT
3yljLpTZjgyI7AXvuXTCQtez5Ix3Xr+6V/h8h5I5J0eVSkdawzgV1tcXdMu+dzcyq+5US6TJRZsH
MWKPLMJfylWFIugfHiyF7M68fe/7XxpFV+NCngpSHBrr7cH87hSKhsxn/JzVE031eZU+PZOzHpc2
j8HYrCqmSijivzTzCcEkFtsnkRnvX8L/jjPX3KdDuhtNUQCZqRkoHlYddp4OIK5+DUmfg3U0m3DJ
05JiIgq1sZWektmQIdmDyUWH2z7J4Op2Q0dfV6B1uprDacmj/sHBEB9O0Tv2w3qM6PAIY+dyxuQp
63wRvbIcF3FpGXGNqj/Kt5vsM8nAI3PkccAoodIJdw+xXKvbKGQg2tZP6+IAP24r29wRRxaRvBKJ
gZbTpSHGBvHwbf7myjG1HPsDq9c0v/Qf4pvvOvZqfaCwm7GcLEzLQZi843UqiAgdNDIgRAtWnv4S
XasJG5Rd+XcN2fj7ShnqCkUVEmKkBTAMroO+BtnjM/OWGdQHSLTys4EzkH8R6kgV8oFiYkECjJ7Y
4v4848MLevAbLekju0tywDmNxhHMQrhPDOmTjMUhwrhPHplWO5hVin2+CknjM53aGRAZd25rQ/Z2
IHwiwfQ0+h6lB8uGBX8j655uUmMOs0zjkm0MQC8IJn+9Hl2vJy0jEdnbMoyyVXvrMXmLSa6wvVpF
lMTIAIVOS0ptDImqjWamRn7grBzXVEdo+pEcFxWuS/DIisAXu6UnB375dc90KJ5cGlwgXve9l8EG
WmJ8TiwEQ92DZAuSaiOPomJLMWJpLIcnU5JG2hCsNf+fMMCfMtveF5xL7qHENR2aSsstk7iuBq0s
CNRdkSJEgYmYHiZ0CjQeJOrnl5AOQuPgEh/3ISFNyajIfaxFWgSHz1eK5ojKsq4+AXCNFbJx+zEr
oXlGoAxgOn8VrzDEd8TNu93WjAWqUNS0UEsAgeh9L4LXgcwZV0912JOFK8d5JkBh30Pu4B4ZB0XW
h0OnJPCVcB/9ZFrkUVFa1ujNA3jZ6Cd4WerusuXifNF6Yl6H3Qmy8WzKFbmuJ8ZQrdmlipPLFhx+
itFAmmL/MGg7y0ISHEx7VJ/pmQvZYKXaMfmPcvZNgDKX2Oy0+qhR9DhNglkobCV4HNekUcErrhzm
8N14Z+rZT+FO2yVxKFvRu2OTTG3115b0mJaBvTXFdn9PrlgHUFndRfRdygrKW/BH1spLzL0fohiH
F6FoxxKglWHn07ctWAz8737wDRAUfGgChsHn07ATEzPK0kQDhkaRiFmTsGg7liRxfvAHVGBwsSgf
NWHc7DlrXGJWtE0CWVX/afKP+0zN6FhVTB1Qb+bluJGjdIPw7jsljCb/fqrRhQa+p0eGNpMQINfF
6r6YlJeQR9im4NO1jsctmHrIiu3WLNoPNfVt9UhXWfkvHFTy3Uj44dWlgUGdRFozTulw+2W5AaKG
6o+qE7lwFmLu22M5VYm8o6WNneWVN8EhZtAP9m7WUv5tR1HdzXKAv89hxEKRJ8Ijvi8UDzLwssYF
akRa3+g51GpsTa6Yby7Y0W1u7M+qTn/DiUFRfNJVcTIvOuYHmX8I3lCSsSWUVsbMfMRweH4CvKCT
tCaGycttvAogaPHY0eAXElK5i0Wbxonzbhv23EOV1w8XbxCf2TIzmKqeRg1/v779Sf/UnRMauftB
kiCZtwMoDOJV0dMv2rc7QlZUiy25y4H3RxgtRu+rs91YR9G8xz53V96JgR1/9SppKgFAElZCuUVB
gXNOHIW9fNny2/nIT7c4QQS1WzIBb3/5gGCiuK50zkcRRCxT/ggm93exHUYjN3ynOAAOZCt3Oobq
RB/cogCK/GtVxQ39qB6cIka43Nt8FZRYJXEjzrPQmI6k+45l+M239XCfMneV2s4dHAhDlCZrENAk
V27UISx19OetNLQA6Pr+AtbYYxgcBhb3Y9KZX4pCltHXyUcqc8j7YR2l56IM0WRwL4K6DOkw0BRm
vvzQYWRMqRn+Db3WpE8MW3gUbdiK7+7YuvN3zE6Zzd0QkExvmkvpBA/HeQoAOum8Y3mA0BKA2Z5/
MPFifVoameVdgGvD/r+YgmIFsNVwEdtwqfUfxIuXJidCGNhKrLNpONkV5q7z5pPRnh2oq0XQDWc7
6SN/i1/7aYw3cQERKvdQs93D7jnLPES9rkYI1GePC7Cxdoni4sMMPhdyWtL3O/MsvHWOO9rwMQY9
KWooaci5+b/9bPfp9VdTtXQdfBlmkzztU18B0oF5j+p4sK9t5J5Wpoq+VhSXbnRS2NmKLJb+BZ4/
56Nad6+RGejRHUgrxGNC8CoJoV1oZp6Yolu4NCcxPKdAlV3z5DJdl2jLV/nj18HUE8psVwTgDe/T
HDFxMBty6vgyLd1kqo08Ad5zzLhGhs4mm5p4TpK2iu+O1X64THSHtmkBFHhFhTtRQxTtArX0q+Gu
5awJDURiAuH7YYsH2s27PDKL9UWSWGkiB6T+Hnf9F5YtPJpiMsDKLKCEcV2P+f6013hSctifIEHG
Z0yv7KS5sPSr2gIk6BSbzjYK4U2qgq0TvkSvhUiVlh+4dkeXDSGcoRkZsevRQ8Cnab7eE+t6wpjC
bjCiW2cRT8kAOonf3fZ60bJr2iex/59+NSqCDOVbxaJHP9jgJviVbewShKJOxuqYe0V6UsPQY0uB
leoaNnXVah7CmMVj/DvcMUQsl5Fv3Z7vMjzlhZWdbRqnicgvWKBEccKALIqMizB2AVOH/qS+iJYv
mrNMqYjuhuendqIDvMQiQAQsUirXEUhbPz/kRwIeUJbySK6tQ5OcvTgJWfHthRvQL0qu10bQ6XQO
1vnI0FbPKW6q+cMxTj8JW0yVxIB8ZP17gQl8/xNSF41IIRaa+YmUWkqsVGoOFNnssOxnLQrPsvhW
5vfnVTbs9oR+/zFG/pj4IN2B5T/4MlPWwQ04CM3e7m0YZpf9NGBJHXzu1n4VH0nyUfI2iP99rxZU
DkQyGZeBL1aMSXiaL3D84CoVXK+FnxZ+PO59ElpdXbEwKcxiIACwxLzfZLyLyhQr42xsZRGYVpOP
abiZHSBV0YpO18wiMh3xR5fgriOsBYS3C8rWiO+UsIG4JoaIYBwLRlreNWWjRrx2trocpXg7zFYB
z6PaubUVF4w+CM9Na5PHgJKooL8Bn8oEC3itgKnWL/jGM8Awj68SZF2LjsmtQ/a1TUiaF+fR+RAL
pRmfB+1eXZpU0QvVUXK+Qu0LEYuqUc+2fkZWPKofQYNK/1iQWgezpUqCBMURfdbBKz5/9UASJdju
UYYFn+H1CWvwZSw2LfaDAmMtdHFTOdPaQcVVMXmjlCGQvnMPhasjb7e4Ntv4mv/RKanS2gIu+d7X
dxQj0py81MgSFlBkIjICEuyzlbLfaJXgJp80thbngG0yVayFVxDDvCmIaVrGDEY+EyV7Bj6K1prn
lDD9dtMC6ucQ7GN1D8yVDsAjB+surRIfTNVyZqRGSbcSBg+vc6CrTGZn0lgk+KjTGl28VEp/ph2f
bDWN1+TAsS2HapnwUZQzcmisUM9q44al2+PFBgyrstKPIMH0bu5/vHk0C8ZomyZ5eh06CV7WTEpN
Az9cMeb2Ok/SNhH9G2ZPYKbjVzzPwnjGeCI9PAgklHUIs0BI2lO/1IJF0ki9Efn+bXo2aa6Er40c
qj/uvov91hSuPQZN/4dgaVCZfxgHAjKZ8s6RS9mJeT4pHU2enDdjatT6piCTE0o+MOsAYZ7uHdox
6orYbT7SFGLlEu+zsMKhsivNoZSSQsbFK8aX11bJKHdIQC/lIWkLMYxKRb6xyuIiXlssv405ym+a
6Y2ikb9i9L253UhPvVOvt4ldl2n5IgkJniRXa6VX7sKRgpEbyA33OhEXqA2cfwG1eHaIHlkDoazI
TVZcf3DnPGBqcAi6Kqck4OvL3nv7xQsIZ26AR7MPK8Hhzf67TSYBsm0I97bikQBj43i2Z+1Uxqx4
/wvoQpYAGkyyUUFPU5QMDhT9WtUcr/epx+PQY9SIoc9OXLrdw/RFaEnPjNLJiCtCHwEnsT8D9B2Y
mqntdSxo1xpf19yHEy4beNSGdphBvU7JEQRYg0u+z6nOrDHBJ/BD0CYSFVKj+6y03AQsrFbgopzm
8qYi72UecQdjm68wd/+r3q+y+V60YqBZsz6PTd+vsTMOdVZVEzNJ3V8poWhfIkGO0Rwwx1RfTf4v
cc4Yd/thP72QEda5nOJtOd/IdQu24PcyKdvDgkkSDV6pEpbNgmi59caGCLVPGYMozPB0NwmzGPzY
W/XZukSJ8qqgZSPgV8wmpdImWpgjZ41LJH6PVSTPF6TEHzmsXs6kh20anAd+KAhoZJZU58zA4fYc
3RK7K3tg04sv3iWxHnwH2l25G9k4WH3E1j+Ty4lVKQE9le31P/JiYyz4W4DUZXAxKg8pdyL/ghLe
fEQVfytpZkRndrthM06qoOruDad7Fi1EQ/rWX0oI3MhydQvIs9gZhQj59GqO45kJHoLGWaB/8rHQ
5vZlgL5rS0yM+2Tl2PUm0s7EVR7JV/eCTY/4aMdECDzboEqY5uTXHWsyq3nofROGprEyE+Z+PQPd
vJCp54sVskaMNu9O+2Y9lM4nPP4aPFUyUd5CUn2bFuV7/sSkC6VumbR42aS2F/MSwcCzam8slTAn
hu7PiJkbj6EH9OE29SEXlTlcEjJxDlQVMUzO14oj+SIVoZCjvvcGWYY8FZm5KvsrjNbYEOn4hs3X
U1tkrVJ8UhGR21rDS5TEFluPmzRu2SeoiS+GIGngSwV9282tBlr2KOU1d/SPZ8Wfz2HaCLEoj3t0
c2CKGP7snh+Uvr5YkApvoiU5SEJWTe8HyowxaveifCVTq5CWKu4azlL3CpZsBnDLe1kqhxU3SisW
5mUksWM7028PeqjO17CbZHLXXDCfHTptY/nM1a93gHPdhHBNMZ5qE8rVZLbkx1IvRZiFM+SUP8U3
P8XBMMaYLIhYyKlrdywbZtkMmFV5HA89/S3+e6hVnsN4PkVsMNCh1wY3GTrHoBmCvCVJ89l3psKK
CbFS8Xj3JSxXJv343pIaW2rOudM/PoPHUbfNGNOMpD92zVsjUEjKTr/R7leJzHN44CqPX4Va1MwZ
YAapcU5T/EW3I+x9UdnBUQXJRtHPdsexajfkKKotY00oTzYYOptY5ehavBTkvj1X+iksQnGGyQje
T4hFMy2dRnIn9kW9hhbR6ajqPmIPbibcOjrmJe8Mi8ytuEZaYgKYaoBMhNY+7rQcXbidnSqozz1l
b7hzZtel4kdlq78xUqRPdZ5NR9nR8ln7I2j9eCiYI2KJ91/zpXO7dE3kJKCQy7WjpHnIPrmt0Z/d
32XIsLN20IgHZW14nvd9YN9RiTEYViJqnNuk52UJzHN9iGKQ1Hjyisy9Jolc7xSRdFuLP+lLi8xD
34Ft384doDnyEiWRgXNjoJAJLYX+Iwkz/UIOKPzGakXlC3pA2gSBfMTr8tez6/K0mk4mj+Zg4guS
9TTcg6Zbjy3TCS6kP8MWgTFsfrqotJ/Uvuwi7gmehYaivW9LngSI0/anXH8vb735MijCwigrZHRc
RKZnE/uyib3aBVksvgEXfnyFnmXaa4DqXcZq+bkZ+k2w2tKuEyfg22Ojx8GFK7lvsS58bgcPfN9s
9nhFp41OVvJurdzd8HlsUG3C3Vzcxomt5JqgY1onbd1ZSWzamj6eRO1agXvHHC1NTsMTZ+K7ExHp
Lm334drZGYVKWRzTyPctTTpD0WZaUgPowmk/sjxOkw8v7SaFCog2LrNYSlajkzpcYEPlH45uXeOG
EjV3Th+1gm0EUnBlBbjZ6VxitE0A32ty5IGr9du5/KqrO94HqbNaeVRMuYqbB73FqTeVxi39XmXR
r2ARZ1PeOuIdIHEHZkx2P6KkBAxxE1twbvaUvkhDv3FRu0TJbQCLlSF2iMPj10xwIl9Ynxy3R45j
cOvFyGQAcSWggJshBFNMHfcZ0/y7UxE9/p4OOA0Zz3dGcLDv0of+s4PztRLqOUNw6EjwF4tKRgXu
O4Hk8a9YYz1lwycR22IXlcY1f4W1AsBCcwbWJiZPhMtl4mLbgR3j/DQyiGeeB/DXNXIsv2BafPvv
jiNgac7HpxEi2zWoF4C70753txK9EUhHZNYnqnzB5X5KI+buKETaF2lpYWTAc7UpyeKpjUl5WIRP
XW3m5fObcU1pHM4fDrwhdBDpo5IjN08VnVficPbD6pDtWsp0LBy13+oZTcCrlOAM4xvWSWEOdqlj
Z1j2GUThFbNM9mHx7qJKYq2I545qGSF+fiQfapA7+GI5GcrDCtnMP88Ij3Zz9vwjuexvjSifVzha
cVhtuNt2kjisnsB7e073Saw89l1yDCUipqKhGt11q6fqubr6mTZIquvi2ewlXZCQU/RTTWgYvJ0O
tR40wUqbE0mndHVb5li6Yswl20gVTl4tohfFBK1YdHc6BTYEiJukSFRuYNNoIIq4UVtf+1CnQZ4j
KYM/WwEVWslPKB9TpGE1nOl1dBVZ94TT1IjPljFrO/LnKvcz++mEyBX/qpzvcHmZerDWtMah/1NW
n5VyPPh3O+iyfHJAHQ6YBri7VsCAn5TIS+GYH09F3XqGcPOkTdwtmiVPYnnHuAke0PefnoPxJL8u
w3lRVjNO09OkwU/Uvwbq+gycVa9LCkPmD7Wzv9YD+GkAxCc0ZUAIDlA7BbyI7AEJFZMo3OmYIcFJ
aoQrXPEd9lLpuVHbVslNibazaJs5bS+qDo1aeTbneHAU7gnIYEzDBh1eecVxEHaMe1vXAQg3WvSD
eSNWoBrEf5RSIQodxfA9YZJkMhYHmObsuwj0gp/VQusFZulEq4rzSrocxd8D3sI5LCEqr59PgsXh
/jIfQhkBM4kUTMy50uCk8tfDWax+1q64EjuD++8Esng2TYu9ycO0uiR9M9W4mJvI07/J0xeoJARK
4bHgr6ZA50eD3bBXrFbxT/ULnUc6hqfHnk+E+frHnHFFZ86CMnomOQb5nwRBJ8hkzDkiLu9N89aX
WyFD/CArRsDv1hE9RR9gU1g2o00DLdXN4m9aW9tSQigSD4F7D0yqw+e7uVqCypLMe5scI0mmX7iE
izVVLHyz5qjZdKYSxIEWF73IYMrs82+6kkW/Z24jxIkFPHuLCq89sNHwyx7XX4RsUgrzqs5DAJzk
M5mQ8oR/Om3jxdHsZuexnPEZFTzMOvsWhGKK0YY1aCmJq+Uzcg10l4JGCqQUyBdreKJeIqJ5BkME
wphBpmHSpOIHUbJZGHOn4dG6UYntdUbXyS2rKcMkyCF3nSktSM8qWaLo7pfZVJRS1Ia9MehGrRzZ
lRWABkEAriFYlVSxbF/B8loEvpxqpLrdG98oWU5htqpQblrPNfOX7NCX41teZpxBuGuYmSQI86FB
ByEVBafcwTXWlvO1JVBRNlhl5vQ8mKND7WQjmgE06cv8KFKjplRR/6sqmTWnWIIrN19snaAQ7Ynb
xw76zgOs21Khdhv2e56fr7rGW+TQp9N8eKuajiVq/I/R3NGKbU4OSGcbEHEy6lP2/Kn8+i+0ED1z
l3KHJ8Nhhz3LPXhPr7Pb2HUI5pS3uS/54s46uA2pJ7NiGxErSIcRLxIaOAhYGkk1kU/ZfR5CSTlW
swdrZf3DoU9kXkoIu/KYVe5zuss32a/m37ttbrXxRu1LXWMFaI25E60C+W4x/nFJ1a7P+rRar3hS
8AOxYzEzNs+AjXXHG8HgCROswybBFelJptmrNSFUYpiB9vq+MwthkgiiG5xVxYCeoxG+N27RKBTX
aVhFsOYn0vwCAcfJQ7GVkFjdh8cVW9b6k+nnSZ58cR8/litNF6UVZLIB5NhnSAbbF+R5yxib+Z4M
RUVevOE8L3ZjUYKOP9Ila7cnolVSvI2NEQ//knUOHywwxBc+bgx/shJqnr8EIiZsX6gMnIYwCSpu
9RnzfWqzlbukZ2p3E+UmXq2L0wWDpykXG80iy/isaUGDJ1eQ2oJJZs3n0Vn7l44GjI9zFyQCyCia
S57t/3k6oDl9hWSAL6cWGmbSTByCoS2X+u3qPccXTYtYRMs1EWvgf2TemDzaA3JxtIQh1Fra6Dn1
9wNhZekpBorfIae4C8qt9UBK5Zqs982tUf+TaRKsIfposzLGrg+oPTFvKw7f/IjuyK+v9BrMOkRU
ir9Kzo4h/ZA0CDNQB1OtUcCuFlN9pa9T+DsLrO7gIqNS7bA5Hzp2IMz/UMf5FLs36cdIJsSqUzCU
mE877T5T+c44oBF9PhrP4j8VlMYFxdNL2zXncPBO9Ga5VLueEUrv2ysIMhlxPFVTEXdtJ3yAyeQU
tyWmEtnICJfi4ag+nEhf/+ndsR/w1V9Yy8gE9CShXq0MlNxVhdHlxmIrm8lw/jdbtSj7+bAvzPoB
z7pNBe3F2qgwRl3WAyu8cTCJC9N6Q8nlDeK2Ts6HsOw63VwdTwIwN3Lz0VdcfxIO4z3NPHBnyKh3
Tf0obcpmIOnH0wbQeHl169ARP1/OpONcL9cmwQugkJUrPiBpSd4jKtkQaGXtvxw5xGZV6Ze7tNbl
xFGKHwUViqXeIxRMSUxgE1IGXMeMmr+wOktrZk89tgj8Y7DFDGVE+X1ZD0PhANSBIAnyemfv8uG2
49ckHe0JEQS+cM2WbuwPMk+UxeVXVXjbFmz3c03/Zwu06Pg9GxuEInbrhWPGsgm45y9o2L0ERnCU
twVxtSpxI9Bs7rxC9VEsK/tzA2GpGgSJuF/ey3mfcRaG929VK6t407KTrWD84aBr1bfCp7BMHuZ9
m/gKDZvp17EjuzwE/y5rNVuHTKDCJ1e6br5hUcTV+cFMC0pTpuk1e/bwpASp3FF/qWQB/Hytk2ZZ
bCUe2Fj51m5adUi7xvwS6DBuhtUnn7mPHXgr21y6mFZYsjiqJ5VOPa+4WMzwUemUnDrHPNroJTkg
xaZMLUTe5Dkhgc5EkI11ZlRdf4ELUGX2lBF6vsnWYEySD6FyNxO4Tx6x6JrNA+OeOV6PIrjjI9MI
C5cyzZxZHuS0Feqrf4vytBSoqXMi84yDgmI9UShK1wjT47wv/iQl7nnPGuU9qGAoG1eQe4pewr6V
FYoMguACP/JuK8+wHXfV5w8PVuNFHZtUmb9wTJQ/mDsettooIs7qneJg3lIM2lItEES7ebJOWZ1S
r86vLABBbvPOkdIg0Sazle7LCboFG0v7CNfE1YSCOHk4NbCDcg/sSCzgZuXxbFxB7jaJsgzBDfDM
VWtMEIyahDoY9O4Gtn9nLhHSkHScytoRcuFpQu5vrzbMNb6ZECrXnTg9IOOnsWHyTlDfEZIOA+MK
tZlGl1mn6WAKrR+4cUycNr+8KyI0ziOnegI7jpV+AR1xSk/mOgetp3JbGxIozKu/woGfwKLxHMPy
3bhUB9GbiaIIv53AOwQt+uuN3B46F2pVD5dhUv4mIG1OkhhslRu1vu55nw0eqOEVDdGsL2V54MO1
D8l18bcqZ/QVO8Rb8Lsjaujg/238/g8fS0bFVfxsNJY7g+Cf+0QK34iAqA53Ry2ZE62YLokAECeb
pkwC2ezNLfTh7M0mUnYfce0l5b8ATKhJuAznMHjDY/i3OxCqOKA7LY+IzUbcKHx9lGJh763d8SLw
w1UGB8g4d/nIS+soSJByKZNKx8+pXaXTztgY5Uag8x7zf/CWy48TV+QriJEnAnxuCxku1m3n5CkE
n/k0p8KofFIvk9RN9o7qfk60qGdO79swxyBg7V8uu2pkYVK/u/aevlsFBivofhD5569uoeEMz+TR
EyNbKS6Gx0gyQ4FVeGlZRFgwDopT71DJ0A9AMFeJA1zjUBQ1/YKZeNyj2Yi/rF+BHLFSCOUVH8o/
/67Yk/TtrLsK66fb1ngY0Kef33ANVnFYTykg+bZNspPDQr+oTRzm+UceCz3NHETre0i5I6F5sf2I
jxVa02je41aH3Fjuxmw5OVQYEZU/tGei7EeiSC8AIrhGie/0iBr4TuPAX5oT8At64vmJ+xNTCoI6
n+OvbC5FMKizzK5SkxRXo3XKSkmyGGKozteiXIBvCfnUACUqxdlI06YXWzoWwHmxE11XF7D/AOyd
636cpkzxLpezFrRnOgAnzBiR82qsgE5nDrCY88MKoqBCByYRNXliCMV6PL0b+PVVgJ+coUvzXmI+
CSrk64/dMCl3Dzrr8vOlbQ5scp/5Rxn4Do7W4nRLLzw8g9wbmm5uFxCY/m0jSePVWvdJd7DmhWFG
f2KaGUE5Csnu2QuHgJ0IlUYj0mX2zb+On8/GDuthnQwPYjBDJXwQzpYml7SjW16D/0s5q0t/uDbF
cG5BG6oNCgoXR0T6M5RnelxG0sGuyPnK9keMn+2UIX/KF7ifhN0zkiEuUSE33HHu9HRyvYOOow20
nnslEbUj2fo1wX6nvRIifpFpvN+MlqRJIb673UPN35tVieDMn2/pVhasq9RUMYFSD7BA8gDT6od9
FmAi0PieYr+XMDIp1u2cfy0NXd1rg4YU/++l9de59EuJmHR0z2znVDmVWotLK+E55euo21ibFex1
m8UHTiSr0RmftQ5HspUPAaJMXRTizAdBLBOcgKAa6gMahoDa2cztldXb7iffZIPk1pnF09KYB6jX
vEDD4em+qudbXWu34O7r0vt2qbwLBsb3WzdG0SjV+5ZnqPlQUQa2om2iKZInLhN643q0D0jBZr8e
l8TidIKxljupRek+nP9DeJxTXk8yB0gDyGJD9GnvXkDNmEQBI9CyPfBrvuFkoyNG4DNEiKLFo7f1
B8HMdDhv44CGwDYaTAbV5LuQShaN0IMDgWTXa2C0I1lsvHbzw14+wKbaa0+zZyPSNE3iFyePa94v
htC6mRH0zjMihl+q2+Lw7RdMH3p5pkiNQFq3knayHg4pIJshsLmnR0WHwWI+m26Phg+1Ji+HF+GI
j/GeoODrmzF9Iar9ipFh9kamqLNs9pKW3cKIWhITub88pyqjY4fjrRvCEUIkLPw67LTq8Zb0EzvR
+x9WxNe4gJbVXnaqTyPq3yleB8d1BkNoHak/IFZdemRJGi10eqnVohE+nSRDmlY9kQZWlqFcw9pp
gRx9rvovtNCCvyWUZgqHEJ2HI2W3ewf6Ts2rFa8sSCmwKq652uJhV/c17huPCNivl5nfpQ4xDLg/
lVmbDJt0JLr47/Ri8hdr38MK3iYkixCdtwJ0pF990hc1aNX2ONfDr7Z8kB6NQkKV0TikeHKLrcG2
clciUoJR0o+XALuv6xYF5uCp5vKGyQDoIQbzvcsa/GeQImwr53VJMaAK8p2D0XexR5crRpqhbI5R
U1qJx81rgM2tc1wHPp/0xRmERaIw4o5NwlMf3TW7iK8K2HQNl++Xq2wFVGrcI4tfVZe6Q+lMKBgZ
hP+o1eNBiK2QKC4QF4HaGi+EYCk4rjb3Lpqiz8oOeGbEt7VP6d3KnO8kE8+vIPSu26VDbu7Bg+6F
SRlUNK/43Q4/qjmjNnrhkBg8yQuRsywI8uidsWef8ZeeS7iola5PQtLPvWtWvhmlyl8MrEIUJfGT
2S+wxFb93SBUyBxnGeto5Dp7cqivN0M2MuXJHscXkbZkH1tCuqpbbQvHWhMjYPGhc5zWzXfzvR2h
Nf+bmdWEPt+X+2O/tqciYIXx2f3rasMaT5adxxz2pZudk09ZDGGjjCyabIowx54jNu4rod3yvmxM
5auE2mqOsMHUgaEr97/ES4wdeOkmu4wfzmJJggNSjFq7af2TIGBIZOWCDc56Xeb91bru2DjpCo5z
fhovammgq/WGu9Tye7Uktym2G1fAUykIv7pB5rpPulflOT0IvdVe8Uxgvq1yQL1/xcgY2Hijm0y3
3aUU7WNvnFr8639RZucjKFxx1qkygP+GSxe/sAmoKV6muMEqa3CkFkp10J3r293dHMzgAAailk7E
c54V5148uMfz2zGAiyTUYo7FRfFEMcnFMPCh/MoK9jV+5CPIm09s6i+P9dlze8Wpb7HCDtOPUmy+
gtB4GTSgql4aK4+jLRDLw+6WBmcOt/9zpf4B15s2aOrcr1QjidHDlCHttgafTYxwVamea6PIox8o
b4wTnWakCuM5nC9mKh8jm8vTyizBEc8KZK1T+Lk2yoCd/b+Sne8V67KCL9Gq99/AtH8H1G/fl7OP
W5WYrcc0QKsjXwndDfvpbWMKDc7dS9DOjUO3GE6QH7soG/MsPd0bOa1sdao460+eyIOsR/luukjM
Ho5ce5/QAApAayZZT/F9dx49hsnHUdmeeNICpvkaONjqNCchYqADWuQMn5IhUm1ExbcK96wO3Ps9
UQ3q/7Huiq+Uqtu4VjT0iX+9D9+6Do33zjEPvdnY2uc5hbo7GmKelsMKuLKRdfqi1d8GTSzqW8eD
3NVSqVYW8ssCD9kvsEy8lq9zLQ5i2Ts9sm4Yh5Snt8d6N1LgLxYOOlU5cvXgX0iiKpeZjVzZijWR
ZA6qdzt4hEOWXKiNqLH8HSZG5g5tPy4PBS3rhkKQZ2sY/R5HtoXivUv6p0n2PQnYIyHCZHvE35nv
HUonKi8SsPVhbRcySfDBrl2bWcRK/JXeuYmGyB9TmHTtbEw5IoYf6uLXaaJyB9NuLQ9rUh7mxXdZ
q1XN+kljgfKR8/TOCgOjIdP82JPwuywes74BK5PAugklAV4QwXJiWOKwodfYk0qmuP9T8mHBPqUE
DCn/jk1wq3sqAnqtbrOT/NZM3FMGJf+Kjf4gLYCFaoDegi5d1iVgjV21MLQU8Wbkih+FwiKAFzg8
hMdSEfyXvZLohpCR4Is3Xmiv53Yot0RKT8xhADX5YLYa/SSk8zQlpkjLsqy5Q3uLAQTfedpaKTPV
UfKIEAeAwrO8eZi9Ti9P2qvD68qDAfyC5xeTnlaSmGcqLNr97DEo/sC9TDTPNgIqEDK3CcJCuPkK
myQvvZmi5TjJ8BI/cUcDIfhTsDd2S7fvHc0Dc27VT1Ja/WnaysONB7IsVa0Hcve3jCkIazl8cr7c
ckO5r6e+s7Ua/oBDhIsDpIVZYjFtYIcU1ZLVEniCxp8UWDE0KBlAxAZYD4n8NPmt4umtG29Utc03
bQih9Gb1QjkHWOD3Z2PgB+qrz7nU1VTyPp1Jx6Y29/N4VSaLl4ck29nkKz5pAVt79eSyuodKuQUN
l0/oa4gc0lk2psoYnk3h169fUm2sV/0aZi4P630t88L1hGc3WSJm3Lj97XBXk/++h5xxNNjeBQdP
L5/WUImniEEhuJguz2yFA7E7izFvBVA3fIVHJOmZqIKDqolVQderiemE6/VoAoy22eaLgRcSgndd
f73faAzwgCDLWWYR4NJjxf5g5RZKQMBgjh1/b+uwMWalO6ZNAYHZAGj0xKFk5ubN8FugGL0oNxxw
tsTGdqG4+smb4wPsLKlFRPTscffRFc2JF5RHoCdIsUKHid4vA/FEwnLuA54uK8xGvOnPXwEglPKc
FCNQWZeIeqwZXxS5xKhflp7R8tuGbs32QXhKqqvH+1Z1VBmpDy+fLKWkFu8pOn/+uUynD83qhB+L
8q0AORqr3wL6YHvWVSm6A4/NzL9I1GEIgqmO5DIbxBh7222leGVEUMG0KAlKTEFiC1mNsLCqWUEv
daCwffoPl8wFaEiUzUpu13XC7zTnwI48OgSSBNepyf9tMOZf6/F5cCShANABdOlCpU3Y0fg5qxSd
Eg1vpW/kmCbMQWd3EmpSkYchf/YBYbzMrSlkwGzbfWuXfKjttYuXLyesxL80gowJNSktiagaErDH
zveiGmBUCzzzCPxC6AtLe9nrPWw+JXlT1Pe4Nc7nU/cC4Zm1lz1uiqIYvDLfHIaGbGrhStDqiaoq
K6i4ZIgFMTI1nOw0/ABUhB7WKxB4dYTEW7c2orzXNowJ5jYDTt6qoNxP5R4t9vtgkiC71CXfaHLG
pdBHlP22bRo9DvC71QOsbGanRP7RIEic64INHQmnczyY+wThhXi5kryH9ScjnJbTk6UAZXAhGsAo
dHhQ/qaVYVIsAWgcgl8NDehGGKsP5bi0ZtBcBid6BCwzphq/g0LfS8vrKxA7yn/prC6kb3zXv4u/
OR351XjgBZAT+9KfnKRorUaUT4XNTTzmPIGeS5tJUUDCAQmo23QMnUYwL1o3Q/+BNeTfRYJ2aHPl
0mOw/Ykj4GfGOBYb3wf0mDKIsd0p8i/tlY/DT32E8GurEKyvzBuX4gbQecZyWZMbhzSPK1vIP7lu
/pg24z7s6ES3J8RzJtjiPSBE1sfswPlwDuQVt6SqtQ18N1Yv+FFv4SfB2cuNu74cW1+hugmT9DN2
PkcaJ1Af6gLiQ56KGXYEKp4ARhidHwtI61bD0zyZxwtK/acbDwts0dVakzhVtOt53wdPK0I3iyIn
E0GFju1Z07jiUYqoOatrjOimLxkoqYur/xyM3BooI+E1KwJFSsRzRq8ViYmtb5WU/VDnUWftk/2Q
CEWzWqzh/ZNpkj/pQpFUb1wVoqnx+BWCmoZhGZ+SBqpQxDtPqgZQQ6bLeBhDJA75LMbuTv9RZ9Ud
H56d7fWPWotT4Ymfms6qhRPa3vhKwYao2KaCQo8XpPeZ0+pmoU5p+QvzJHBh4nS8g7H5lXJXRF/A
1kl7gxgJj4Q3onWESJYOHP2jgBNoyqEfvMM7/KN02A0diyrHGexXHPCP9AfnoeY9V0ZVMV+KhAf7
zdYDymyjPGIXi3XnMrSL6o0oiiZxA8+wFk02h+LI32kqcghbD6qn3lVQqNbkDA0oiQAjGgx3WrTx
mCld2D5uEIpBQ3uHrbGz6EyKKI7sCkC9PIgEzlkmOH8Sokju8BHnf5vlc5vsjOIiw2oj9uqspCx4
CCWWs/AzlvfgtI0c8Ei0mY47Y7Uk+UsOUTNZTZPa+Odi9GQCYNIKB4z5fyDu4UMCBoX3bNPg2ImQ
aIUQ7na8kI1s3O3/l3bCys6XSNEwFDu/WRYSaXSUN2x+DKTOEsULnJsGAcwlsaLzn6mpfphmYNjt
srLMCRoNfNXYzg/xErUVIRxJqRNvKRhbwhbFDLbuBCpRClzXCJeXz73hipPACa7A9XtSaJhfw+pQ
TtkRsO6vhi83T3gHC1rFtbLANKFOfNpPKivyTXe4skq6TmFkgEfLtDZKOGctwsOPRnqCK5oH5OaT
bs/u1zdPhgojzwP78bqjvOxlQevhxjhWnEQu3kcLvEpml7Wv/nUhI26IykVYSyPuh2xw6St31x5X
c3my6hH8LHc4Nz2st03mhqg3UpnyDJGfSGuC6ytLwWiLu24cfNkwPd3TAH2iUPxsahb1+vN45W2T
E6oBMrOjiSnjfNvw979t7Q6cV3dY8xwjdorg8CVeWce699279R8K/MrsQLHcXHJYJYRG2P8pSjih
zARiYeatoz+o31MFOz/kd6ZDjBTrSelOLBtLQStLgZc3SMVBA8Me2IgIzVdbApXWHQibFtuwXUM3
yriImtc+/bQhoXaT86OZfpX5V+89zVh+OAMhSDSpKEKmJ4Bf0Gi7jO6LjFqcy+gnVKk3+PUmPDP1
RQWOYp80/60AfMHhH2iTue5MueyxbcvJbY55iFJ0EDo/hT5niyetLiUThcY7Ck+fGQEmXlHNoF41
ZyCDctZX7PWWuf+xXfQZFY/yDux8kIY7+MDyI35kQeKgkXCkvjB5XH3evBM9skyfTja0QIRTXbR3
4Wyx5eiy0aYsbYXli6ydCcTodHaQL24EVWqF2lbOPFA4vC5GspCPgbbEbjl5eMVTPzwlUB6w+El7
/+CK+NT2/8TVIpo+djaCUkU9qLA6fhIT6c0ZkU4LFcszv6PsJ5rFvL33xLVtkM4aXgTprp0LbY6D
EdxaH52PtxsUxJRxafCklANBFZKgImsVvRjoBEynYkNTCgCQIkpmEOcOIZyH0GeBeR2jkMBSK7nW
iN5FmIzIvnfgdqc8BefiC+bROX+p2c4kglnZljCzKHuvkBZ8mWfAgUJRPcoPh3j9mbfz+VdKhAXL
rOxssw/7wIp1VfqyeV03L9NNcm14rHIH91JdG8qNRAG8i2adGrTo+050520NbQZa7k+WgUGji5g/
z86M2yzf3gSF4B5RMp6xdno+E/2NF+RaB7wd+ml1kWDGKSUwRydo3l99Hr9Ar4raNHYnLHg1siAF
CFsBbYrjuJsrjCdm2Caf0QahIytI5krTJdhilThmWQ7OfMhCd1hSGASSC6/7FFHNVdDvtMD/uaCy
ru03OtvSmMw8aoCf0Bu1941tMbVqW2otv2/QtjNBofM1pBJT/VksCx69mLiZHkH1vFjb9nUftlva
SGVgnSozMbog/Hjp6FqUhMQ1tZa09RsWbFFDO8v29IrR0fMjwXJVAyUK5qihlbbHb8Yx7C/ld/OR
eYnUeDC/ygkLbtl6CGv8Vq8hooZ9VlEuYAPA39d862T0ssXqEuyvpcthsMDAVhVTPR8+ygVRdhkB
DqkKoLZz3XKkkCVEX/W5BThy0yYyLv5FdtZFujY2/XjA4SCfHk+aGg3As8lPHm5h3hiKFsgw/niM
oBVaFNnk//9sXFQ1Empr5YbyK3PXZbmwV9lWk42RJJOGZk8LJTaG3q9s43bQkUkBNAqkPX+AovAa
Fd1k1MSdK5Fv90u+QS3wr3YuPwVl71xKP8/bVFxZNvAOT55V8lwRkhoP/yflNWQYndYuU3z+VEuz
iLFMzAbGkLyUUSnHfQ4GgoHmLjPNtJ4OFqTub8/YTN+FR6SMKa2PiIKbspl0V2TywpC4TAXflbyY
Ek28gMrpRsuiYus4xmJitXBhVwwtM39GNNKyCa1q98a2Zk8/XJxfVlBaI3WK4o5Housbny2DfDN3
UZZVrbKY1dOTAKHFb0bRFw5myLY5CCl2INsfL39CxrKSy95pkP2EPlKrEzoIZGhUkghWLAPRIOLj
+yDNcFF9YCvPs05a6a4g/EPAXXq/AgiZQtARdoBqoRxWDpoA4Qa5fhAkY6pan9+V44B2MA8dOBa8
X+uE45bO/m3CsMnlnqlqldel+M4SpC36oCJ3z24ye95rECpqt+m6/oK2gLCL90L9hHPxs+wHVzNQ
5a766dzGlLQBscqT/pWbiXnHS+9z5n9pfBe2qP8ItbADhwNdZjjqztA8bLrWoW6OfnaCqgSY8c4c
9H8lExyyadULsviAC5G4moaIaw0O7aGMKICyz9TD0NpNdD6lLq/LhqWriWduuD3JDIiZWGHeA+gi
a6KoMi1MC/+p2yYk/5QGBm8rvbNGIyRxYDej1Y0s7EVXukQbb8LEW1n61rf8rlJY7cX6teKmOqvS
2yi/CQF6xseQw8XS4rYiE3KT9WBXiCDsvWXCgDMbHHssqpe3XsS8tfCjAagIttKFA1PHv47KGJjG
WxazrzFP0aGHLrBplda4PC0sfjGsY5WyLQxDG894HhCgtu45jdvk+yeK5YGFC/um1bhFyEIMMQ+/
rtU8ztRl3HuNPi2qaDWpbI67rknt+3CgzeGBfOd/bxPIgqNqGMCm6aFHhNkKwk41gO4jQ2UKIh79
RRW3dV+RRBO0CBYzzw9uNloPuIQJnULzqGGj2wc25fr2J7HJn01G/En3hBc8sBjAvhL4RShtJkIj
w2jQ+wEshYNB5EW7aJvWxVeho8qNPdwPVuIF6s+7n6FniMqAs9/pj1flnlVYyeTUnhdDFK/9U588
Y4D0Qv+tOiMlAZG0k8z0rw1NhXz/DoSzzanGl5FOZBqSors1zbVYmP//ndgkpBn25IbvVpfm0AWh
eaJg2Q6EZ12o0i0j5vMEP+hflXUK/VuKrkKb4+TNdVZJiQAXSVwbvvwjS6TaUe4JVlQNn2QHlflQ
RHAquwvtFzG5uNZfx9+oMXQ6tPmO5DSm6x/G+8lE+Dr/tJSMJIauBstCpTqNUywA+5iE4MpjXamJ
xYw2CglB8JWItegZt6fEvGbLCwkkw4d9pqKaMjI6FWr5mo1Uf3bmFT+TZR2z2alTjfcIXnXlZSEV
rO2PPM/jnZrym+BqfiyDupsxyzcQXHuQExQRMhdYD2uDoX+yfz6qEcjUAkf+edP+p562Rw0/QpvO
YkAUaZz08u0I3hLZVCEXuLDFk/Yp3wug70kPfEgqOLqizqDjTqw7wZMTJ7JsY//JSlLsF8pPC5EA
uWSsC0xXROQsBHTSq3DY6VQyZ7YODxG5NmjGy1eJDnjXNG8KDsE+A/tjn+AjQLseuSwV/vnAnUzD
lx9ncPqVbWp6L/RTEkdQ1y252HSJNbfqI4XEy3uHlXtg5U2QRN1q9YEOHU/u/0t2BMAiIx3P074Q
QeTbB1k3m/5wKqitzZZQnXBijesnbqLAgc1UpyXhHj9oEWaz0CqSSD9mO2HY8Stgl/a08k/CdBbX
D4xKOTJakcQu6NepNCYKpUs5Y2DoMk2HjsOjB5aiaPraDA8TRRbi3EyD44/sPzL185Rnf2q1bDmt
DN0PKxx4JC/7mDpeaWqzRx2eH6+L/WwJDbAvoVOQ+T+nO/JxmgE0eFxZpn5Kl1MSt5yXQFNWrSbw
Y/QSrcFjE5fo2QdH2TDaNbTip24bWffQY6u1lclXB1RB7mRIdY5FlSlsYpbexB16/3vvVyM76YvI
TyVtgNw8Gv3L1GXpkM9yCWcIN4PDiWyDYB+VFOw5WBD1Ic7uCQ/ijCKDzIFtkyFtnbq1mSZMLNFk
0yIbQDaYk7DnDIk5igShoyxWJsXq4tjdZJguiS+DeyrHaSbZL11FL2tUGgiP6+KWS1HFnIxI8vNK
HzuZM0gH1r3AxeyEft+Bh5FJ/farlraB3T1ZYueAR0Cq8tLWbmjm6GyEty1rDDtZBhZi3iQu5wzb
Jn62IdrQLS/0XpQS5n2K5tNjX39+okujFbI6TeX2SHRyejvbn8XKOGO07MmAYVg53NQufqSCzJuZ
JP56iMdYlSe/ZrtsbO0b8J8WWNttp3u+SDN+FV3DEtMDFmIEV07B/a5CWVpF/++/wU3PMRQ/7PT7
rU8DU22W+1UPOWzac3Aw9Ct3R7dUd4MUbHdm3fk2y45kl0pYXLoxDVj2ZujEjhPX1hAH6En9HWM7
TE+8buh8IQq0mxJhuqTYvErhHvH94hEhXeZaA8nbnmuJUEPxsWBaHR8yfVJitlegtzb7L9YhHMUx
uycv9P48RRRXgYQ1W/IumZa08tIXIoLthYFIKfCBZWDsVO32DenP19n97Ud4aHCCEqkiwW+BV6f9
+lKCfpSgP3YrHJWAw5j5NCIAgdLofVfkw8eaxRc6dVBv9CWnR2qSBkUEakdnqGgt04ojBlU2XEsI
XPp3q99CHnqfhGR5jTKJk4+JGFnjanDrogWansbNO5EqEpUUIrnURQX12nPCmMfzcNzVIAxRSxqm
4RViknSx03iFOafzbwDr+8iONn2cW8eMCbXb4fnI+P0B95Zp9oADTakiEAS+zWxPKDSQYLZLmP+/
8JovN8ryt7VG/DyvS4847JGHwxtEb4aSy01KJ2Y05TYOYDoPFb4uU8scYsmPEt3/sdV+9l7Gssxb
RESM3YcQUVsznQyL/0CtZy4aUz0Bn7nx5J141C4uMl0qO4AU2hO5xNX/bOUibsPB8uHyjL6mamFE
lr/GTuExwFMxgJuLF6tGDGk5snWBAZ08RdRGY7lPPzp4Dn6mmEyjSYXDLkxmD/Q/11QUDNp+lG8s
37hgvxo5gojiafmwXc4Jet0hcP6h/osGyVCYHQBGCKhCuEaw3aLitTYWhGU/zUPyUbgRwJ8Tf/Sa
eYwR4K7ONfgeSBx1U1Dcs2aBOrKwui/K/gomYdzXb7garZXngL4iThbeci2Fi2/Ouxla6gXGdhuP
7/q7RvaMBeTcS2SGUDFw3p9eMRtKPfnwEqGYwgSLoVNF4deNdpD0XJVEdtEIkm1sWjG/PSkKYQTu
805+Wtp7MOdAHLQcEH/N5iRxikpdYBKlQ5RDx4I/rwk4WIcdpkiGCnheyh278xY7L+DQNzc6Ul9o
txT13JQ+udKIA2hrDF6xIY/1nsj6sOvcYapGkT1DLEc0Eb/wHs+sdFINXSd5/E9N+Qh7XfIVKErM
wqwXLjStFrzfv2/9iP/xaRl2OnDDMPuUnDkS5nn5nn7xoF6aXg1vtrpJAEpPQ1dw/sVncDTF95lx
65879CgAliZWBr8671p+4UYZRzAnUWInC2pC+ZjUqkArVWZ0VJDsEeS3S4rTHXdaTzkdt5AIOzUv
TuhXzc437CCjueMM9XIYfOFnp7sr4c84tzSJMpal9T1I4d1wYn28VPrw+gwWr3DZeOVb2WspEnSl
cJn4iVpk2teTD/AwfN8UcMz8E6bWJPTySGBSyAil1MJN/qJOIzpy4V11Fm8eAyqjvi4BGDBCl1CB
oFSRa7RSYXfSMlskNke63TwPrfKh4F4AxoHLYtueL6anKV+lGDUoPqvdUv+V/VGAiG3o5XDX2fcI
sMDPzMFK4MqsNVuA9w4OoiG7I6hw8ccaO5eK5HVsfye6g2NH/5ORi/GrUQXBXSgEGyEsku3jKW51
OsdfiTrG7VgttWTmElADBTDCI8ux4iHItgllKBfv7t9hbl/7c/T1oiKrnEh9gE70OM8elnKJgHGt
aP+EIRSIkGjY4GzQJt1l2M9d9dDs2ohA4Wtz5t2fc/1HOYgQCZwBYiHtxWhfXlBmxMv+RViU8lB7
elfmNDMFi5bTqsZbFjTsNcTwtpre7Pdog1yonbPiOe0lw0ZDQn6Yf1rwxYMm4Rmh8yxNgtuB+bMM
azIPckvwXYRuXS8qHI1T6hjNPwLqpECml/FDRw9yJr83iBvelYPt2d31G7jfZ8B7SxFfkGQzzoSA
5DVcwtPS1h/dU7SIgLLldyxI9SihMWroPUYZ13ucc3n3TdSnv3pcoYcQzlWvgiFD6ec2weJfKWkx
EkI8QZhbE++7phmzNRh2/fTyAxDeRUH5FrxSWjJcifphG3QoDR6lVcosUPApSFTCXdmG2Fjs+rSX
leKM/iIzKrFjY/EPRo357k6jmCr3UEQvjmC//1eSGMm6u1kw1ZxP7ca0tfhAkGxc1lftfviVORMu
OVBp0QM070TmRI8l7acdBBUxevDGtD2CRbgZnt1oO00yhXfb6cfWmX1HNE1TjCOoRSm9nffggdFb
Q2dxxyofkyI5GJQn2yYmB7AnPQyM0xgfv26G2I3VRxeokKCNIoDdUykdnQPaFOYMXbAVbPZWl3ZD
tdp6ZQzqhIpXjRGv13gsOUW/EXxTGkqPudFdjD7Qsiy0e9LPoYDHqIiBvW/ZpB0PpBP9brDEWZ+q
O3u+IKb8QMT+Jt4xjhsl3/JpqEZKGPL/DpMJwuitIfj1jbPofGcc7qL+v7wIEJU8ZMXNM4d6YbZS
DDF/ACFNjkBvUsy8VXGvewSTTpbLLYXs/aUvkinu3mAwo0RXc5Iv8UFKOdriw8WOJCQl5gccrk9U
88l0aGbfuYU/cQnGd9z8IfmfiOupyJmgc2qEOOYdE79/Qu6lWA9ij+/r2EAULREauqntrgO4Bx2o
0SmQ2pzU09d8XW+v/jBHaN+cagbFEc8xVMkCQjj8bd07yP7pQcWcnRJGlcNvv6LzEorcTM2yOmeD
gMODClOT3UV4oklzSzrOSbMh/4vxsMAOe8CPJOM+B2oCwIUphZ0ruc41no7hlsRIQo6Sy4zpCUqh
oD38xmovYIgBjbWEN/UBsQBwrCAowgHV8JH54sWMGxOH+EOp3Fi+pEftOn+YN0Rc8SOZdp602V/f
qIF+9TSAPGAO10v87KLM0rVytWx7E+iO20jDYK2Vwj1ga3FG4n/XurZ33nj3G5gwesf5YzuOW/KJ
3qKDiUOdmpC5n9+6htWdYHG1FZOmA7aQEZo8KKrNvrIP9kQxA8xLM8Xxz+AIDfFHEe4Uugjy4YgH
EPupIbATAyhJ5jHmJIYz1IzYuKaDbYdy+gbzX8n/vO2vMEs7PJGIulsZmW9vEaxmYzYJDeDdBNHq
rLrgH2WTVRhNkximuhQ99+j7A9kEDrV9Ne77wUXl04Pa9/aLqIGzNR2X6C0+eLyIeildYfeiaolH
TCYzi3p3lRORS/V+EqdiI2qJMKZ8dmKoirXEReraAmoO9zd7rYTimtLUA1ciU727J/3XjzbYpPs5
ZygtfMOu3OvpM++Pmgy6YY7uVmmTUr9JJSJKFlcP9w2ZGOfIGv8l2mlOW+GipNpxOXHWHchMr6wo
AIQhixtlUDxv5S2T7k9fK3viX0B1lAChI6G46htIcsukC1yzX4AukawF3/CwWf1pvwz6iZjS4gE5
iQ/ziR4w9K+5gy8zzCsjBcbnFo2Vz6ImXNrosOl1e3WVGv1Fk17JsY71SXvD3JboQPnWAhEUyN61
pU7Y9Gkkqlhik35TCXF+b61CU5NZ6snNz7gHjBmqFMbMzT15iCYKY6TWoHtPNVxw1AQHpeUDd6hk
rRo4XCvfAU8vWU7b4eCiwAZDZQb7HPtQX+3b23HC8+JJCzDu2wSD+h8N7GK65ej73A+44fmqEAKR
wuLRs0Nn1+gCM67dsof2mR53YmKoQGPQGx13CimQ+Q4tLvWgNEx189EwNL0bbn1ZTUGdOX4OCX4t
j94otdUhocILBOP6T9fKpiJkcnYK8pqWzM0uzoZkYOHSzmly9relDW9HD5vpPH1xXI6OHlMzWZNF
BG4YGCCCpR4HhozfPr49KYI2iA+nnxL+8KEN+A7doX1rOekzD5xEB4Co/tOLEWg9CfcmolDNSv1y
HcdZygXJAHoM2yngCYUAlT4zrxF45X+l4+RRrNavZwyaW25sXdpl2gayMKYgC8NKjEgyUJ7/dMUK
B8ZWDDG0wEfOs3PMu/j+aAXloNTcEQsS6LMVmIFiiEMzwbfw3TZ4kyBtnflKLiqEXOTFvE+TlRjq
U5r4YtE8TARC5UgdAwigy5mC86m+sLTBRed7/19gXY5qw4zWyDmyzWjBSexFigawQsiqpK17TnCF
Ff4Up9Rq4pcIssVwwsmnWwMfpKhMi2LuAU09N5hDHiBQQzUyekbBuB9xTSEiYk1q7w2OW1IHSe+W
HtreDzc+hEbM016SHalSoqvWYUldHVJbJ283iIKs6Zi6FCl+q2/XBuAwlRkRxMjkIXk64iekXBId
88EFIIlD+bLjzCoVlj3t+EhVi70sPSmZb+vkl7IqnQM/C5bArTuHH0CphmA3Sz/spo6aG/oXFRIN
FMdDXDBrD+Rl5F+Crjdzh3mtaEBl+lrJlUKtWhmxdVcRQh3k7ANzXhUqyi+RMrejdLOldrHqgwlR
RVX60BEVK5Fvm/pfZ+l2flzi3MKNXnCtBBUpVKXBYwduVolBtR3ekL49z3EARkJFFWU3KpMo5CqV
bvjiX1YwGWEKly8Sz452asRYz8JPziWlxcGwlE7KeZDC2zx9RixBFYzK0dG7QvRDiti0/z3MyvrL
dUycWno1VYw8nBY6uUTjdIZXX2R7Z5rpDoDqNh/FnFtjPIMR+0CzbRo+kDcgNNbOWHOQROGH1UGB
nYikl7Lnp4/RnpApHfO5x75+tsv4ye/FyJ7oUulLhHTp7hYZR1qm1m7BnRDRQCMba7fxuBySe7jj
lG6dbgM3i/cbJu2O6+yl2DyYFGvP5Z8TyU4YpuxgO3bofRbhCVUnTAzFDphxZyk7USnHsfHDDdO9
YCqQZ0YMgNoCc+tzNjdKYGfYh8covQVnV6Z5jgVsUcUpDiLVsEkWmNmJoSBwT18sHm5bDEd9H8Dd
rsyY7YA5GFbbNHssApl9TYJasa2DTpI2ZEZRA7dN0Y0nR856+gwqstkMprqQPaBQeFCencr4ejQC
2LifcGm4zXGFE75KyGr5+jLmufMpuJ3Li0W/olQKp1llCAt+z27b6ek+KHHg6k2yPnrXq8uY26yT
YZhR/OkZK0EqfF0xZ1QN2EpdvqUqnkT5lahNpP0SEe0cLptOYGwPZ0xgQjHcHCYVgTn3XRvaFRBC
LXI2sboVIfbWukkXSMQLVOAb93oc2ApbVulu4HDZIgG36GXkUIZMCdXtzR2rs0NCBSrhCYUiWkoc
FkDbWz3SjmYfmLgmvCNY9LPl2632GFewEjJO98r02hgwtiOIQ66hlQvLfykdxlv4rX01uMLq9ymM
jnBpt6Qg2vj879Cs3LqzdWohWCUkDB7/aFMRdWRdXqcO33NPyLthc3bzvciR7NRm4qGq23XOgh0g
uxxhwWJzuYSU0hPlvXFG39TvS7bqD65eqO9vwiy4SWMrdTUP4m0QlTw1i+VAKmxjmP2mOVTH/OLG
0PV+q3SMMuhA+sX318viNpc3yiIMPDH8N6AyJ2btK1lpNo77iQ1h6J7PQ81FAJqIVlkHAmYmbWpq
KGTaf4An+dya7MKB8LkzPtMeHQ49MEONfRIJYjK+sLjkiMuSp/fekpBipw1DbJDR5WYDe7o+Jw0C
OH54ejiXXHwPsgCzCElN0L1uFae0hEQZ9m8KxhV6gaCMb5CDjSpRGu9AYrI+NEn1Coda3wII/tGA
HO2v1djNkAhsCKENgsdb/NlmtOhUjwbajZz6f/2qwi+DEteUmd/rmnfd96QYqz4YwUrsrhMEv+QS
oZ7i1c253WrjbMWw/KTZvDFUvHLv7yabHhf6n72wr8Jqzna1M52i+FVHkJHcOSE60zaFL0Yhuktf
mIrrk5DkdsXVLJ/kVIAza8+xdzfl7xDQRN5Oyz/iWQ9HCCMWw1iHLwdL/rsDdcotuY0TIbBN3Z62
2nCKr/byCvGoRF+V23ePl7XfZeA6fbqGAwkwj+lzsYZ6H1sdPDP81oONIIa51tyDMhHbFzQwNRGD
tllwZmZPl66JgbW9kky2rYgBv8zJc0YkbIbm3s7rzcA8/+0f5ZkQfHG+TuRbtVNsu5PpxIGjOcGX
crY0qsmTAKSYkkNJlCvB/x/mCD8vw4gjCf/ZUBC15nZmlKNWTl2Wn30BFTHpc67tuL/4XKVejZKB
SJBEXWCqpRprPPW0jS6ozyHTQXWpZHaxGJDOzH1QM7SEwm2yqc1fHq5SwAn+ajB7D94xZlen5n2T
3zUUvpP29dha37xON61hi77m1VnxCm3EjtqgXj7gOI2Uy5iXR1YXdr0macJ8flFycXDZPMLeWAZL
u+6C6ptyxHNpGdWZbui/KeKWqCgcmeysVzgDeKiJ+E3PEyznQNDzDlGPPpFlbvviNdl3eOyb8g5w
ZH5jw67n7gBYrMqS8PiOVxu9zSPUtbjNCZMxb9jfKbnW7o5L7q+jA7oke7tEAVCz7MwlcHkdCI8V
FS3xpZZg/ckGuJRWSlic9U3ZDmI8DlVmLUZYxy0tpXUOmpj5gHsxjMeUC+L7UGeW5EDPFRC2AzpS
Ocv2/AjMZxCeu5En+fgCtQYCe4GSnPkCkDrP9K1ZwCwBJKuUeOQJtHTRIBv5yb4uUgx3/MvTsZhE
hxWAT8CRUXyOTJ0IZ678g5C7qZ0NkJ0mgoodROLWRutALpKBmduEMR1YDqcfdJopkTJUgYIVlsOa
d+uggocWqnoR0o/RKa2NQ3LfYYkCKNgCbCogEcKleyCE2U3bi8WLHrW/EYY5/xEYiptvxeqRUtQf
0gBhMlxtFtpRC+ofHKzkdV3Bb6GRlssDl92XcFt+zI01dpfYdGAQglqRk4OD3CyHQEd83K0NdieC
Sn0fICy9v/FNI/FZAIDgk/rJScqmwA3Y6Y4mDsCTw75FEBRGo2jrPlnrlrtnxLtT2bC92H0GrhUL
Dvmz5caiRUJaelpSrj1XY3JesUdzzzLlsXpv/NXAVgCQkao30LyX7tmaVLYpKtbFw7sg4C1hPcFb
NUORMb3Sf/QILZhvF78SDfAcUf/OkYrB9KxRSO3UyM+Nw7BWeeGQROUV1D1YDlfB7Dox8y5b3a01
0W80RU+BJ1sNg2mI6afDzZFnovRcE7NkAFO3iken5+Xsmsd9sqkbwDJZBymrYryT3dU1QpnJjWQD
jjR6164AKJ3px5E81N+Q8KakJNzqD+whduye1wwXJkysX8TgPgYgBJeRiSaUsltAJQG/Vo+sYBE+
mqivjDd1xwf3EQ6e0umoi93ib82JK4d++xAXzgjouhWA1oTmWLUbeNFkkSnhEVRfeuIeh0NofeR3
k0haVsAfEgeha71Oj1jXPth0DI4Y7eE20MAVoZyDrD+WNPThGcJ/ZfLZLI3H/ixg4afUcOdCYS2N
LyWLVhBMfz1BjVSZlcHNx7WM7ioOvGFp+xt/VgsCI4K4prvEcgcdVtyd7vlsIysih08FyhE5ahmA
/P7KosLUEybXd1SbRHYt5/sc246g6a2MUZwdAWcMy5YPuIP5IY12xy5b0BwzfJwXkfdzS7yJJyFs
wTGJIBBix5KLgRfot7sILEVdLRgVzyXdJa0ILeQ0n5OJKItTcgr7w+SfYgHsHwUpnmvBvBMa77M+
OtDuF49AXIGZcTuW0VDdFhmo5vdeFcVzhcujPsuUZZFZiFIk3MZl6ojO8Ae/capIhbJrd+gSmjpa
2mSiv4J2DXCN9d7u5t/yaXzUkM/t74XU3c36xyUrJroqm/BukdIlwB7ouoXjbeK/oTI5tLtbUvRL
tp4VE80ly7kVNq1f2xckUGtNpHY3w2ufj6mnRqNb+lQhWfMOLgCkTH4GqDA31I/SCOvQzs7qw9xP
f2J/WakVWrISsj4My3Co7Gxo5EVNVF4Mbpka3RIKRHydyvhdbPoQzoTQUjKXyC+Ph5NDrpnVIoqf
MK8RjB/xE+vH6wXGbLs/flQbmrPXfmOtBlVm2ZWXlDasvQWamKOZNw/4HNQitiI/zy7CYPXukA3X
WpM3t3ljJJNPWRm+D+aNkH3zcBHQ57J+sBEwN0IvUd7XtV3aOO3ylJ9at4FgmJ2u7FV2qVLz+qNd
KyCNIEotZeDYP0P1kcXUEILxvKcJyNQGo/BNUQnXMs34DkpQBJaKWup1eFXnGHpxNtKqKh+wel4Z
mQ5UbLh7HqKJ5x7y5TrckJSk80YgZNOeFDZBp8jHMV2pDgjR3t2IUY0lADPapNO+WuTcAhc27Kfq
x9W0G32B9ZlKYRNm6OsqdAEC2gujxaFOhXxFbohl21fAXbYAPqqbN79Fl+Ss2IiUFMHd5zXJAE17
MDqBT6PpJYX8y2pFTAqFlZeY6FkjynagJ3N9rxFLh5eaY76Z6MohO0cNzAtdwsShgUQr0wcUuRgX
8wKgE+PXEU0/BkQKbSyTHT6NU+GidrOM6ZL7QUbUIf/9WCpyl1qkm+JS4cx8+axFA5TntuUflYrq
9lMdKMoldpAR/kI8i0UtmnYwzp6e8wLoz9yvVFb3/wXG4bSpLTEhaDUSfKjp4MN7S2tHb/fWu6d9
g442abUa7YFJM8kOin3soYg7V+IRX6RHjqHin4+tUqDQ3PgVPS9E+rfeSIo5wdfGHcPQFpbON+D6
/QGQCPZE47VYnDg35MHYwRPyoxM+X4pPUIenizS9BgrS0hceJXYc0Gd7raWpCGMVSuZLE9wnXp4f
XgUS9Z+jO/9dgw6hWDlpaDKt3vF35E9hzZmGl6yFJqdXB9ovYA3S4+xPeaLYAiK1RyKew4YmLJUT
NBTHvuGwt5s7R3DvoEi+TsRcSm3SS+q5J51PrdC/LPS63Au0QQPZVRAYqbZHnYaMu07fvSdHV9Cu
LgKenWsChpqsyASiBEpFBnXCmO6nLeN/zYZvNNKg3e5HQBU4dbSvWOr8J7vZE8LBEfCDy2CUUFRR
+rJ1SoH1H7lLB3uGVk7zQj3WXumEblrJXOAb73I5UID+Abvq9/0aKxTYdQ4XKc+J2rVvR7Q3hD9m
g3cZk5z2youVabk0Ng8p2hVU39Pc1NXgAkfNoeH1TeycH5VV/CKh2mzZmOMj+CU/odfz9rAhJIC+
zeBCm8LSGWTCP7PUnIYyYTpV4OU6fk9Gs5QK+7K4HmsSaq+Du0u6Y8syBap351l/BR9KRegYEFbW
d7Cnb/uUnLgKccEiXJ9jpR8xgI6giyO3EygtJYGcgPmHgAEhVM/ekrUZ1oJ1D2DxLK9eEpgDPFUD
Je7qpv9x8rNRSUFAHpUuGeQm6hzJi+V9bVB+/iiDiLQvwrGlhlYN2xhrScw3KBagI0tgCrXNph92
Ku0DBBxcUeuheZvK0Pnru+/Ydxg30grk64cQgPEXyTuXuLE40lQhlzyxtyHjJ2/mbyE0TJWAaub6
1LVQ14bYVYQT9gtz+Nxe2sUtol9LZYZcu4FftgwbwoqKnkRx5GdUUVCrHXSWkUgIg0HAMOAIq8OO
TIniqQzpCjz+q/0X6SFl359gmANlQL5qlmTrkGJ+tv8ZAMH18qFJB8lWBNpn2Aff1OGybmpR7JrQ
GZhY7/O5bRvyWI4yeqR7n1sj58v5+B+f3Ce5/JyShM73s1Ft/GSDFU0njHx5fZBCZiFogB9rfb5H
TC502zTbFORcjcSZ7f89NHhOwIgyAa0/7O4en7Nhm+xhsw/QZHpOJ70cCmF2rdiK4q8B9wSXKA1e
KtKLEx82Jxur54X8emAlordXXLY3qzrf/BltB7S5TK0QLVW2aO0tW7oRFOcNus5eRqyzaaqX9CcF
TRosISai4Q9Q6X5lPmqCOEJIkhYDU+vBL9w0GhXJXG9PZc1Sc4RxXR7N0iGBZV3b+MUNo7UoMJrO
qSFNdblD7j50Bq60sEhGVjveW+lIbeJ066N6PzWKoGYdYnqMbbpbNcW85IEXWiA3S5D0aSSBqnmB
RfvoN6mcmBnqvUX0/6MeamWpOaScjNrGBS0VWVeRX5PC+CovYGx8N+4wgvCUCFsjT0pFBYRHkR8i
wPds9LsFAtDp+6INBYbkjKQFHGdx6Te8DzAOOkSrQhZnxzsjtqQZMh5MCXzKkXXEWMwpqucT6KKH
tNni70hV/jqNotMd31eLi1sQiohCat2sY083+REx+RZI9cAttKd1CNueaC0WSiBmoskgl6pGujP4
YyMOjCFJ8suDytMSjD3IoeGctIt+bZX2j/EHl5I/JVUxvXATLhXDimT9vbNxhpd07TR5ECh1lNG6
CWozGpAYgv/9cV/PIjGVAb8ajYZJoMb85bco42Dmgycba8lFaEm3WrQBS+qhugsLP5FFrYtKcU8J
TwCyRpDbKj331fAdbMaqakd1gztWZUniz0Q6KMQA8zMYv8Ik9m7iOd646s/YF3nm84bYVmlbwmN8
Je7LlhjRWJn5gGm3lQHah77icgRKxExdgsN6+8tMWLE0+NF+lH47TXQYRj/HKYuqFQntZdxMTaR3
5KQI1YzjmR6MJEki4uYQZLRA9PVJILJPiSmuvd4dhsCR6KmUYGoDZNtP/DbvQqrWRq77/RidFIbz
lmOpzh3ImIP7GiKkLkqVAr2fOV5KjB/e7ZT54qze98IwAJqd4fCwBAH2wmVs3h8C1QEn+tt+sbJ4
w3VD3ZCW8u5jpLsKIxabRcuwngcy+KJ3jLHdP1ZOb2/88f9ooKerx+ArhoWQcP6genNsLiZBRiIH
dnh9u3KKnbYlE/dmMfc1XUURn1Hu4QRI2Vw/x3/qmUF62yDg0yNEM8MS63bdQmsQr/sbZimyuKCi
KkTsbCq+XCKbfGvYQekdj8HiYHBasr6QbG3LdGmNIIX3j9k4lt8CcFVoZRkonkOWUOxYTX9Om7i8
DGB7aghdJuDQSzoju/xXf76Jc25qghbOGqbIKmYpPyviPygZWjAQ/yp6pGl4zVZDPx93QDR8wZTj
Pt+XdNmgk5PGSZh+A8b1T/lspHnDLQzl1bB9wSg2ZzbC7+bNTE94wLqidI2i34JjrCQudbDWMgHp
5KUcpcvB5R5kKVBYbYTJq5Sb6ceUh6brjzoVx2wVtY4g8Az23EXg/Q81/TDYlX8vfBuE3JoZZ7t4
TFz0gwOrLddrQY3yssV70dE7Om501KE4zeWaC0p08sh1uebGpPQJ01ShbSLel+8BQHpJF8MEVm5x
YWz3pwPpZbCoaLzpZY4IrJv1dM5kdpYVzr/dKF5O3n3ElmgFL+V9HwR5Igap4o8OJk/reZWDeeh4
1sUw2O19oZFZpDiRsRwZv3FsNCmdOYXhtiIefeZF1+PpZ4nAicvBe+IWSJsD62oN8A5S8S8SpL60
xLVhVdoOeMLDuAPG/HMEKWcRNoOlZMpfuh1WvqThquRzLkdjKDzcMBGTB09uigWjVyMJWhRlpu0I
6cbs7FZizqgcc2kv4i/n6NAzM2GPsq/Ol56m/ztKsMnGHsEelJPNdn8uxZTBoz4+3J2atWX/Jf/5
wn5lYJwBSK60rez5ZZhqGzq73daFYzAX2YQAmXkzWXXFIFCfqHtajlkwzT79YjQEJaDNJLjwi86v
JydAGuHkifbFfyKLEC7FGPYY0MH+odLdR46yn5gprCKlUo1G7pIqOaE/HnkMWyjnDnaqijN7wLw+
Xh6le0vNZrB1rvlHmcwohh93wajxwyTW9RdnVsT/0zi20x/e/VgNQI4xcUGs9rZslypSH6H+gtAb
spnyv+5o+1c76Pq1E33D1gGYSLBixvPa/4d8tSZ54Y0m2XuB17HLQPgeoMrphTIlyWnNs3IkGnON
uLaenvBLI/49sbwnY5Q+942TYBxV0FSxrYTOWhsj270aKYSQrxuiDV798lZfvJGWl3c0A7g5VVuX
kLIktghKIiUxxL1fT4rZSus93KP5Y/L8yh396kdTqmMbA6JxIjwOyzGUTGf1qXufWcx81uR9kU/R
/xMf4nYXHYtrdKx2X+SvPSMY9KRbmTt31FtDVVDT9h0w4+r7ytU87d62CZ5YdLJI1M4RfmIZHlL9
YX5Z2DYyj3FFsDNMTciDm3QoifSSbG08p5Pw63hxgCJwOSBglUpWjGiw4DHk6wxQRCRwUED2Qqev
gL7v3HNix5t9b82DvgXQbIEeBmJJma8p6dFo1a6F+jM0EyAVoB9mmfLGwa9117R2y2gX52s7HXnI
H3JIYehPC2bfPNoQ7i6HLysG4/8SCgmfffSHFQN6Z7hpwTRsUFM4MqjhD0WCqn+SeZCQbrmacqvE
39TNOknAKP718N8g1oEzD6+XMOc78LdueZFINVvC0pWGsHWI2Cgzs5Jgh88YTCIrOmZg49l8Keq2
Xh8TXrk1VWnjJjkUjsDBsQJEZ2I2x1jXwiJqtK/VMEdRqqCH86eIBmGXmdN9FZlKZLKqJ8IrRpwD
GOXqiAI4OkKYZwXabq1y6t9CYCkKDZ6VgX3NMxQtHKuEz9Zd07JXkS2C2w6gVOucq5YA9emzFOm4
fGFBVLXg45uVw/YlHGUNJgI5IChjagi7lxkUlczbhHx8UcT+Gpkz/DGWC5kTOxQ7AgAUU48o32qk
bKfVONS6PdBFJo4wVE9k5SXLoGvsPUNKQ+UUM5ZDdB9eQDwMEv5ADmss3d3cKtENc3M6iwtLoHbL
SnWprQdX1DnqdQxYfBa1hsyjSa4RmHhml+2lXR62a+K6bhXVSuzyuhAdxgnc4XyeDNeQWN2mJ+Xr
NSjfkx783Xb2flbZlc3wEZgRDoi1xiBPczlQeM4dLqATsNcAA8aMNPY27ZoKBNustO43Ry7A6pXs
3H26sHQt4Ei/kj0M2ojg9QgqjLB4LBVr1yOMmRQQuEIBzugWPkc4wQq/27/U3wTPIgDbSiT+kL4q
KI6EeHmOqqkVO48cXBLwCrDP/dKH+ANl/+Lw8pmCQkMAcaQdx5iKO4nkFxN0btFXUJUYO1uuj8Z9
2UrY6KiiOQmT769KOIM7kAU4ILiuedc0lvKFihbbZNa4Ne0PwO/BqWB+MzwcCa9j8KpJiuslG+BO
IfGB8yevjqrVb74E5jTw/BzE8GOqlv00ZWlm5GC+ULSk+EPySpuWBPjJ0cXX8DkLLUcGjf3UMWQa
N1rdu6gQcNGAxoi5BKPI3C3YPAENj5iVQqC9GcAE8xFsww6PQy4EE5srPbghd1i8eJjXhEtueb1J
U/p+cVyN3EroAgVLNeWRnhor4bEYrqDkd+E1sUUG46DpVfjQxoOgB3DCmwEGtvnfAOx9J+Gg2Y2S
EA0qYtxNjR4Yei7GzotK4uMH4KTnhIKY/CIptOddM5IWzh7X7uOfzTRU5nLSs6si0SJfym6Tz4mL
tY5GhqdxHr8r+oJiv3Yr3J9q6Rlhd6k7NbyvmPMq3wjYB7iQK38n2Tlo7slTKLMRRu7CtLDVH8lR
eNRqqXqwPzEcvsiYVerswLcD5A9+gKCdEG4lCHkX7Zyt7PGM6PW0SARhz6ZPP1FHsY6qBpG7yuW6
Wuxmx33tpZA2w2FDmIGygfdIBOSnwucPN1yn0riklDmuII67EoZH0b22StL5Gtvn+fFyxwsopg/j
4ikFIfpaaoQUs9R3T0QeA4roT5eOj2HeeK4SEX369RP6kRTPva2UApRllVT4gvyn5u+azfzxksGB
marMPaSHpPCxJtBQDAqWNRYC4Cfr8k7I9n7QH02OiOaXoTXLivsfKtPOa4w/+BxLPKf4qTMI2Mzv
qaN3h0UgsCtCmGkSU7ojl4zo3AsgVMoKE08RqfqqPvCpYSk8GiHWyO4O9T74Otu1lRjLTKdUAUcL
9TeMCsO8GYP9D1ZQzuVVwoO9e/fHoiJPkAcy/UjpdWo5aD+1qQ2djmR02jWRRbuoaND0z/256uhP
wtNfmPHRfhyCFtvCrNI4eHOuvT7a4JyOnbOKcWxJ4T5NgERpQCu05TOjJVUsfqPDM9pcJ6UXgSLx
4oTtgoZsd6OuoEI3uGc+sycdR+z/hJaYC4d/wOX122lO5VhCQ5MbZtwJrYOqSHsFtfANx2qfkJwt
i8SmntYZWtRvvRwdYvJJ7K3a3oZoO9yqFTK7TrbHhcUNffQw4nTXTP9bsUnyIWkiB4p59ef7AU9u
n+J+6waXNJ8jGF/6eyLDwPqyPmJykvxm+CBU1l05DYIimgVOQU8Jo7cBJxOMt/qSlDIIZxyMd1dd
cTZSMD8zMYcJCOVc+cfzXMwkXvQigveaXhJG33VCzBzDVqmaYNWDRaKP989FmBByR4FG9ZiofLlt
Kj1NRLMCilZde1gSz5iClNe0Rqjt12cOBMLqu7mXYJgJ0y+inVc3zVy89Gi3R2EfcnwjfNp3yjNk
3QzRdy+AUD14Z0UGTUU/j0xfAklz9Z5HscyHThXHdkRNSNmZwjSu4L99uJKSDKXZoGPjLVgOzV+2
HIQ2tmMWF3XKLaYC2AC1HDV06E5FyVh9M459/8tPYPB4cnQjov6Y+s6j95C5F93rCcfguLtcc9Di
erSuBcMQwurTOoU/CKdLfMBywOnbwu7DhKg/jlu48IU7qNJa4mIZjoH9qd8HB1cvHDQBajENL4SW
ULHsinaB+7hxjPUmAmypoXcS0zlYH7pHJFug/SU+DryTeizbfQWtXeEYa21+SySzffJrWLa0B5LQ
D4LkcGuNRh9cbpgkoXVrHcezkUjDL+gqouOZEHrkbbivRo0tCcyijKSJQd1ChmYkRC/WxCgVRu6F
RF5Mp6wsxY0bbwNsYDO8XMNdJS8POVGWoWtbL4U/RhcbCjHKdirnRigpaHXtJkC8JHZ0tIJ4gBs5
B1/07p4cA239koU8WZErZKzHALcYaIMkRTHN8i4OCJCN5zcZc8bDO5iYSAPaIDMFpXtjH9qRNgfR
cZ1ZJz3rV+RvWCNV6kCkZrHz75/SZDDlo9J1Rf8hxH4PMNSiibXRgo/bgPETCVyVzMKJCx+3KUOr
HqVrKJhSvEqbM9EMzlTH5jW7hK92RpNIwDnv+bQ/z4CfOoKnU53WvpPnET5tX4BGGZUo/1rQ79KC
HeFnWZL1Os0lghlCwgzoOwzoS8eFCH0ZPdf67Q/22KvAsxun1xxnGxZJiVCx/c/jGO+mzifXvYDQ
hTOKhxqTEk6n/lyutsJsFDgu79L3ASINPG988EDc9EAg46Bdz7Nle8K+aBlbYKHVTyfCgjMmmMEo
ugtNUGfUPi2dIFeJOl9JLuqxsWUvsmotGWx9CgHAi62osKkWAA1nsNPcxnUVDcN4LErfBs3FbigV
QWemz56132km8XtXA4XOjEJ67JNGSmOQSja0n7NIH8VZn20DsDwZfpp7X/ssHDdDlKPh2SxJeNs0
m1mHxeba0p67oQL6pGC7OsUhx2oWddvcz8CGkanVxNz/BbbdcvI9LZ2mnoh1jxACUmttqTH1EPjU
s5uBEEFz8HCGyBtX6It/DXtoF9uoX0oIQ/fK9G1diC9AvhLHNr/XXk3x7UC9dHD90eNmxRNjkU6j
6Rnv9xaIZXUJTnwoB7cxhx2bFHDWl4j57RNVf56M+YAQJ+aXEMIoJQ0JC/ZZGcoDNm8iCwv07OUB
roh61hUNIg5sB3OyZ1AcJ4WHb7iHYrTiveBrve61bgDlj8w0wPEkANlPfOMMAuZaOgOMLllap5Nh
7kIqDQ9F0J5gHSCzkDjHVw+2EsCGGTA8A5TyhyX39e0xE3oxBHrzcljIUKyMKoz4EJEUrYVmDaP0
FR0zBDnAvt9EjXsy3ROdaJxM2Cez8w02mdnNqJdghGtyNpUyJ0haVPdrXmXAxLMzsnQtgn9nHI6d
ayy+d4oWFd5Ibp3RDXbLgnLAkdUssDnPuXLz/vwnX4u9JBZL/Ax+lupG2ZY8jXROslTueup4Tm2N
DMF5XkquqTEs5AOeuqfMEOjrRbbRkJ6OVzp+sQMgj7YB4S2SLl7B968MhDHKhC/nbLT+oulqdrNp
ppEuA/LndWTzWL7L+4jSym4l0DZCSzGW5sY1BLbwArh1XkjuC6VJqbjfRhNA+U/qLcUaXGBiFkV8
QjoUa9kjL/W/7Arue7xJ8E606tDcWQUrU9Le5LCsdjRvDywzqJq4drRmcLCanXDUUUORdcz/DGix
L3ag2RnW3Y0FsCHuLrBHPHMZi/BbeuAXV7m4kz4cPuLhOkiTcvq4E20iGYmK+9VRMK6kWLfSMk3K
9t+WfD3i2tN0Vo9v0d6C6F/+WgtehVsVykWcxG9WwRhK8qQPmM08AGT4BP94BKQ5NXWrbDdHIA4e
er5xOZb1jr56oXI3uESbq2bb3vcf4k+vu2q5t8KTJjR+Rq3wB61/Ud4P6a8aL/vx1iuemmGWab0U
2Dt6bYWkoN//SM0tau3XiYfLJhbVskV3sEI5vzBwKbxUQKrjzKoah1Ttw2IjBNUZI1xPzCrqbxke
HDWUQJX3tKjPnQscDtQ7P2clfSqBjZx3FQ6fh5sV0n4XeBf15o/n9ilP6x4Cz61nljQXoEQJbBUx
WccXuwyKfavmNnHT4EMeXGmLzLnZPSVfD3I5/5Nmeu6g0roxs0rn+pAIbXTcG598ZcwNQJfzTosX
vlHAyuzApf8OGneAEFDnTlpCImODCU8K6MWYtgIKMSaUpxT9SgkCRluBm/814uSBc2F+VZhn+VBx
bJtW9bhDXV/RhUeU96VrK1VaSZZ39m0UcdEVMROd7D03xE9//n9Bb/KgUM95GRW8js8lUI3pfSNC
SqC+/3a77wZ3EQTyPf38awLMyPQGJoLkxa4WugT2/anWivz6VOWtEZcs5WgHNqRqWRISoH5qThd/
odujzYRJArVb4wyrRCWvg9QuD5oiV1WLMXzfo45tOFCGtxcB4wRgyE0XT3DzYL6MV2FxUTUjvgQl
JV5GFmZC92nPV/1H4FH7aajWW+OaKahn9LSdZd24VN0CaNYCCvworM3ocgdzvGpgGmDC5sr9YLz7
ydbn5sPTK8rjm8FJPvrPMkQTV5o5ncafhYOx8qXeHJWvAxDP43Pxvv+bkPzrh6UeEoygwm8DpXZX
bQbyESe540wu5mfYp/WG3L9G5Uv2KaqX8xaPDrGHYwSbiUmZ4NlMmRii6SL0/HfvHPrFZ36I1Hhe
zQc0RO2IHlr+MfW7Sn14P2IUnuYSWwQH2+oA589/gd/DKx3oprvcKo/w6d/GvF+9WOq2Z6PHivY6
YkT7e0lsHDYls9Kz76elvVcElRpbr6yGEyNjj2m4PQ8drTuY/fL3XO1CSY+Qnkgd0l3ppAbZ7exS
IOCJq0I9DIIa6uqJby78JJsvXagnsGSJOZEcZse5Ey+lHTOQ3FOTfJSh0RFgiwkDOSFIc37IAS/e
BzU85A0BqzMLks8vJABw7A9LyKGwtmbk8nyfl1FS+9zbaq8YxGkGf0qgbbJhAgywbcMe6mMD26wF
ZXIU56mXnP03lXC3759eYt8m6NN6vbC8qwDaOFLoM4Vqk3J3yNyMNcXHSGwh6xMfNdA79hZroLkb
dIEMZDo6+tQA76BTlDOGsa4Z4s1bzmkaZYcXMbnxlyGBvgbY3Yr2fmMCRuCSO4IN3r982Zz7xjgR
fUA4yDjz0razRUYucv4GKPfr3Bajs/SVNAD0kCWmYlnqaVa4FT9/QkS2+9bUVjd2FRxwX9PLzOjD
Kb6I/qG8VO6Ap3W0Y4PMB4arL1L15I60gITsaaIIf3xmHsoVZqAa/OOenj4i+czyqzj3ldyAeHab
D2ekqpcq9BTdw83hSMovZeUgrpco723bnzTPvp9ejPmVJ3v0u82mKAc4vTki4tbDxXSq6HSfTxfw
v4mlq2IJ8AOK3kj3lfuuA64XmkvELbbiwEuHcYvGGAsRa/7EIuZK260tdxQovAXBw82xPWgTrUeg
FmP8CgzEzbCrOzhy9wy7Yzm/s9LQ4O8wHuN5ftKiGnqpgfiBwOTmSqrycuVZ2hnqXcVBxgXzjhnY
4CTSFQ0n4fwJIKuMSb+z8Lgqm1CGYjq/I+xvNnkBD8fMPvdk59ODGgAlxr/aKQBZ1j/dd/5FwWTL
bLZqF0YUioCsyjtEK8ShJm4yi/c/cx4cOCcWORC/YvgcSN1QKMoB/MWWZQE9c51VlMCRU4dKCC4l
NAf47uwCDpmp0K2uxQ/snjCvdxwB1L2WoqFkFmxJ9L/KcpsGz0n+bu2eX6ySeMLEtpC/U0RGiRnB
rko30s3k/4yd5cxlTrcy6SoLfSnnHL3qUJlb0UfDHYpixfOzl8pkq8zfUIc1bdABaadCleGvH7i7
DoGqcOHatjq/MHJoFxPzvDaEitJ9kYZtMg7WBq5jEFcaYkWtu1OfEs9bK4yWG+t9fvgiVasSDi68
nV4ohROaZFc3YS1/bDImI5LkTPFve3a7MDlfJKmFWlAxoCYgXQoShe4z8fW5GtQNKdQr4rkaqFhq
FXXb6DIMzA1XRo6QxZPTU0fMHAY6f7mA6LX89QRBdOYomMjOIrxtaF13DBsX95/LxrPCVlF2kBa6
ZWK5w+wF0Em3xf5HVFrPFcDHE4rsI78ay2JiL51lS1qg4QcWc27D2vjYFAFDAa5xGm3n3f4jdYYR
jzmnIewqO2LBqXKa63eusP6Jd0MLMrDXp+KBrkNzEgOlydsnja1+cSCA7xfsJrditVogTUFaKF8n
wmQig9xCXS8OK1XT25WUXr0GGWcFAC38sraYMVqz0bJHZau9UPsSEWuaMIKjyu0s9yQqYvFFtUCv
+d4UmQ+LXH6siqXNzqnvb7a7isIJH6aqgM0ZBs6HMCOJvfmFbclO7PSABJrh+SZCLrN6sGQmW1xV
z6hQ/AtUNBo/op8+8OUoWvpGSI3Z+NmeuBX89MaPeaJ8awXRRVrAw5SEY9VGL7jlkw53PA7eyhdw
EnZWedmjVj1KtIyxhw/RZpw+lY4C6h4tC8D1kou+ldGQOCD4BLuq9L20pbM/Gyg5H4DCgqUxvNXa
Jdz6bGpesgP3WsNvyxvcnNKTbGEULvIKw+dRSTk6pmlLnKzB3aiYwkvD6I0Yh/X+dJ9/8+Z7rHyP
q2tFOITLkEy81i4vA6Irb7CcoroOhiO0rGZb9B6KOEIT8QIJuuQIvGKmDmZbuTE9bnB/qh2/HE3K
1mS6K8u1xj0NDXcyXQrp9+FPoUc5sGiR8DNDlkenwdo1lvFGQYP5AsXB3zvYtHM29LZPXMShmd2O
HV4sDl1bi7jcCuYFvyRDXahHkh8Tua0Drqp+S1neRA/bGhD4FCinL1T9g/Pmm910N9lES+0zhdZQ
Uj83JjqyVqDfTIMq05J463qUgoPc4Jk40jCGFBm68OTfkWLyPs52z6dfnU8VDdjuqnhf1mycwzRF
Olf4Hv/zY+cXYBIULe+w6G+mg03KBRhkkvO4J42mrIU+36Le5RglC2EAZbvjOJFrVGaAggPBszZJ
uynMnboj7HAkHHM60n/NuxJkEhHA5O3y7GCFeDQUA2qQlnSmO+KSzoTLiry2XlJvPj0/xHMsgLaM
aED5xt8XnezF0wXJxGt21Lk4jIAPg8wknvqbEusrexMsX8qE7BR/8o3vGwY14+Ct3BntemU7kHWV
QIarw9N1+lMyU9BhXHQSOnizNasE0qzocX4XtToTH2nqMJLY3l/Dh1mh0UY8uDsQwHyCxzPlKqDT
mxy0UV/FUF+ZEDZFfKILRVoB98R+CwX/dcQ6fP99w1n4OFJKxJjj/F2LiXTF7d6DB4lJV6ctkHPa
AIsUoK7FPg4vtyfW6ProHL6VEVUkNSq9hSvwPLTsi9a+PpTRYVSbFrMheX7t4FHDqoQAqY4jLAzk
O+WYEjWdV0gCvXFLMaaCbPyY7Q9xk9H4hEX+ZPsrQ2KgFBzHHhSMYlFLayzIifDTvBeKT4u0wIoY
Dkjehe+0k16pDxLTtbxyaf6V6GHnuNoUlVAFXCzT3q9f1pOPmMFzINq5Y0r4iZFvehKw/Cr0WdAI
XzUgte8CwV1lHOR75byTM+A9aoAVjMzXNSK5yYEq/YTjwsO+tSZr4p3R4VpSJvcrrXhmusN2H3G+
S0oYQuPYSr1sjH0CnYxsyyOVSNlBFcRHBdbt1H/CLlvkioBhEVrl+FNCSqsS4MaSporGKD38lBwO
+QDUqkdJQZjonfHrMqginkfcM0T9l8gmBTRCpUKNwU7RxIceXzCHiJgTy+XU8LPuRGD/v6ElwoTJ
zkuykzTkPsxQv0tKDl9XWzhvDYBgWeHBIR0BKPFi95i5+M+gKbog0HpD4YpwbsdDlNodO0+HrA3G
/kN3zfV3Pa9rcjnXcdc1MriA/PuXmSRi7a4EjTV8rd327y1GiT9WSa3JpsOKE9qJzKWqbtC/YamH
V9Lt+JWKh2rl//aBhMzRHWx/LRTRse75CGhiaYAkXcUHq1RkF4JGtT02Z03t4fVzFGDtAOB5CGOa
h5WDAfRn0B4RD7w1DT0E5MMGfgkx6JYGz2lyAb+KU7ni0Rgt5x0kXXgn2Bs5uyQYF6ognrCJ+wkn
yyvsjh+9mpWF6z4swbke4rpU3B24sOA4k7VNMn8PlgZJnCYJk3T665am7C4W6jZUdYDNHNegiQne
wAO5RwcryTnzlDPYI/+8jHlVDlourdBK9rP/vN7mfpXBAji2NN07D/LgY4dj2uZKCU5FkRjSLWqq
ElUfoVzKBI5QYtzOcyJ7SP0hS7Ucoujk0z2bgN8Y2mO9TvZRe9Po/GB2odV3WepZ6ewMEaSwT2LE
4/ACYXcd0cSmHXC33Ez0Fzv1CmWSzepDRiTbbc0NFX8qwWSyAEpjPPTiQDYaaWVcLXUl9vPey1pZ
yxAMjVaWJIJd0cIVem5ixYnIB5G1NFAfEA8hZzKtlDCH8rQrJWoyRlu5F7lkJ/RkOxr3Nbn5/eBV
e3G9nbdjVXWPH8I6q/MszObxlKlvIxAQub758CZMcWpxOnJTzJG3p3SmwPH8ui1EPe3h9iwNvMcF
f0KL55CCns8A3f8Q6Tfpfa4ylECNAAFjK/RXhfpvqjY9YZjkuQk1KCo2r/qOJqjN8SJ+Sg29t9Qv
+kQPSzhHGZvRujvTIqRFvxD2X4qM+IyRG0V1wxezQpZLHTFWnC0SCcBWF+CJKMMgA+OQjWgIdHGt
FeW/jDPqzJYmO5kmIrGeekn+peIbSSKV8lki3HI9pQBvQOalWG2y1h0gsIMoI/jzbBVO+dblrAfk
ieJaJvGYLss5OwSIcSsP/YxOL9jlVFnuLAyqcR6jUrKy2z2qyShjP29H6VXtkIslqBoam8ePd6j1
DbWZkO6N01skohTiyFMCSSfETNQ9qnOw3TEk0GTE1FU4ADyEO5XU2EZuZ6pv8Gke9VUTXt3myQeG
/+Knal4wi/E+k6xyjSOTSEI0ws3FA7nTqvD/pzEP7nq2waLsIBI1yl5rsa+s/rlOUa2Pta7Lko85
P83AAVzOuFahy08gLKmE/DP4UpOs6r1I7yZA8K0QX0/2Ti/XXvXLdgWlcCj817otbNq3BPiLNKIU
YG85xP9LDxEWcZcKkSlQoB3LOx3+FQin/EE9Qvk1q0Hg/dB+4M9PTskGsjpOaCXagHjqHMMcKGgq
pa4SP4vrbjlXm8TSC0jvFu2VHZ/NIOKgrTbkmTbWxLPvdCCIrv2mzoPcJkOMfgOmMn53uaDnLRtm
YvSF9wv627OyAfLqcziESmUyeOAOOs+YhOUso4eiQc1ynkzNOG26UK9bmHA5/kHszPNfLRT909Km
On27envUot+S9ig/FIDxQopX2Fhairmby7izFYvcQdTq893lgsZR0vnonYioPa50oOzSr9aZPEVp
ob5WHjSDSlZ1bdpXQvYj8rpXibcJPMZuAcWIYWO7ZhnRbLAvcMWYYej1FVwF4t9eGgxgjillpoY8
WU0nGyUjnKRL8BUdhK6h7GrPYc32rR6RlnNGEkMTQxNVgEHljF11K9z/35FecixppfVWabDY9pSu
AeEUz4yiwpr1FoOE3DhJrvC7WwC6D6TW3ojQYlks3JW2GP1E41XIstrRiVgCYx2EHxiU9t2UnTT+
K4QV0WVLkIZhQomjiywxSRbL3BQNnSxIcztmpwapdyEHxXi97zdnuIo1aHJo0eoyHDXGt6NXzaeb
ii+ys4/3jdkWZwyjVUAT3TUP2k+T+gUDj6FScufVa4Twoj6lX9bHogaxIBeR1OFLU2woImByEWYL
4RpuySCOlSHQ2TG/bIAz/or/yxt56Hrbv87Lf6KE9VZlnWV20zAsbfAhYepdESpZzg28YnlqkjRm
XDEA2teIcRYSiQHkUQRPCvHIs4LbgenTKxoGi8zE+uOEnY9JAFyWLpwZ6Iwz/SwvK0hapbD6Y9Ct
PC6PJlErdp14/1/nfIdgiZhfThVgu18Gm1L3pL++aUIl9i/Wsu3GnSOYEpu5L2CAcgi+U6LwEKg9
4tFsjCcEG1OszgVuVAZwKZOCuBgnMzy8lDX1vi0QhG576YFiBXZ25tRUiJSMf8Wv399MtflHG9Hy
rQPaQWfOm7bTVCvxAidD/FyHBNNaQ2B/UzZ83CnwP7BPAdPf/5tgkNuti0N77HOtFD3hfBJVMEnX
+AQn654HUdHb/N7WtjwZtdVZQMMzUcnRSNFYlDYDo1ga0O41TDIlglSpXp8UY/JW6sgFJ4vW+G13
EeMtOD2N64BPflYwi7y15IV5PrlikcUT7j4nTdNgXjHLnCt+wtFC02aSq0oulDG4HqjBUvhJtoG2
aCYxXaTW3TS8ujiQJUmO/5CYrhuXHKqPqrQCQpuX9Wne+UzAzTn7qaPj2PIbGo6JejEfZFetFpWq
II4uw81KFQV+Bdtz0P6SJXZAALcPtwJlKthDFeGXp5dEM5m8OV8vyQdFN81GN0si3P1TcRGVCUVw
SRY4DZpSAjBGmaA2XzZ5oG784LCr+qOP8ppTmNBUaec1n6gVujTwtlFnwjGFUPojHbxp47H1iK4l
o91xIAuOAs8siLfbQdi9tIb1txYf40Jamp4lOucNHZvwl3VtTma+k8n7ilxZR78VyNWtrCHvCfs1
IEd/d8Dfl4vg9U/y08rQ28qvlD+zt1OeUyVLNWvxc/ZWKs75kvZdSOjXxsVf0D6BwMuy6zle0LT7
vF6kdeDpbqBAs3KKOifyUgFezQRBhilXkqSp54+A7AypxsMlVoZP5aIyML1GSij1fNHvAtqGYtYJ
1AzP2GDGWj7ryjNHf4pBfEiaa81PKyz8g1Bgrva72VtmbCTQvoU9gkR3rnSROvgG/wGDa7d5zahK
gcI90hTpj1FZMYKcvrku63keDXS02urppE/VmR/w17nid167hoMutyp4BSyvdHhbEbFJ/UGT87vv
cQxz7BLIzOH4W7Q/BycjAEJDPVNRwRAJyEcz5hAJTNy41ToGlbmXBdIligXBeWfHFsLSNYdhy95n
AEOi++QzlhTOIxvIKrII75N/svimiysw55v6PSiuywgD4OQykbRrn7FCnb631khd4dIRZP8b2b9Z
4V9VnQYgwca2nPVW2J62Gy2wNFEntTo6i7Ige9tvJI12r97LsI8SxfCtrWev1DJ9sMHYBhCdKDWX
wPLHNWALfFBbpATx8Bl50x3C+fb2K1h9UQTBC2y1hfFaoHsbnyJNbfgUfUUckuQxAEqBdBnT9jZf
PqX9SniP/0LPDtUzmvnbKLAPkUjp71p6twerYfkwqCB7U3I41jcIyN48P3Yy8VZE5XL9TF13CASL
x+uoTp8EzB+vIbegLGpmaHXRQ0OHf6djXT9gjWYTm5+2CAdjgGqQ0HwVIVVuGJcGII+hukHLJYmK
I/v5zYcU4ZBNhiyRx2N91D43g7Lr0zNxi/azimIyW9iN6HHURFOL8Ackswce25VAbF/dtH8U4iNx
yo0KFyIFvtH5EC59onpDodIe4uEDITQqMzp0hIWtx+7ZDI0rquaIcltLM+hwWXJSL0uA0u44vPKW
MNiP/Sp0GhNHwDDbOkPfBk6sDtyuMvDC/ZR32d2hGjNWsjs+jfcTTdCpR1Eb1Ko6vl0BygRhHm77
fkJCgcKUHKv5MasWFPDkcif56BDatK3wq9tgQr9Z7lzT0MnkHPzjDoptSy0Da8wXt0YIFKG/YPvH
FJmyPu/94bT5PRIqil1A/AdAu9XFZw8q49nLAMo+NMbPn032JIbE3JV+/TVx3gGHyVTWFQ7z76ZK
/TG402aLfjuY3VlwIXyhP4t6lAf4VIaIORbpyzj74j5hJabMDv6pFBkXbpBGm22/eCYmHbDri9C7
jzwogWhU/UMpFukzIRGnfEVtMoxgEY8YtCk25LdFE8qNuTKV/pf6eTeltOpHJ6ONR1qYoAbKfJvs
CvuMX8wIkl3jQot99xIfHhGX8VfvJHiqdn8hq4+syXFXPOQCGrUzsJW90pT1Zke0rhw1Mrp3+HMI
5l67vhNlxSn+18XO8/U6CDM6f1XEfhKd3YkB0ZF2ePPMYiKAQ+5R4Cmz0gaYdAEj9VlvcJa4pa2b
3mxS/r4ZBd0kgrC9UMePEXSXwy4wJwIuLbVq315n1T9Izb9lGiZMHE61/4pv6SV0TIg7Y2dnOG0C
ObDtE2IY7xYdIwvBUjqCSLZKprzLtHcyuTqjPDMRHMoSk2jDJ9vvOyIemrKutHUYYqvItDDJ3i/+
OXie/Mg/hwJPjMgrqmvUl07uUm0UXC0b3GruLF47m92vDJ8Nxk0fePaYq6FcENNjig4t1rlo91at
GolJVU8xdxWiyaCG2AS/+XuUVNv+gb6mJt7RL4f5KodP8roDCcRhykRRHy/u7pEA6PuFgi5+rKtG
s2tukXEubkUt/TxYOkjxcrmxSJa8Q8VgIhEDQC3QDMWJjfLu0aHmLSr5JaW4s/dl4ODXbw+KQGYo
IGFVQflDXYKFdyRqT/C2NSqvTEJQlSfS/Rw+pwwjiTuvMAQJ43UADw/Lo4nCYdX657e9Ovbq3EZT
v5Z3K7o3Tk3AzQjcOZr6V7yYDYG3mw8wVnuniOOsDIm5zAW2umBECop6rfiwu4/gh8VLzHFHExXA
st2FsquTTIf6pbnDniwsw2cleQf+psTz3NxXuSBfCb+ReW0kZ1WzZbKdomiqM/sEW7LhbNvvZRep
CHDbGIndWjWgCJmbjzXA5WZPUzmRQK1lgRkuT8dwXENEAfSknzPaXxfN+o+RPszKiAxLU9sckKDp
1Kqk0v6ABTSLKliD74ZH58A5WGTFdiqYCsraQuMBKnh3D8nHF2Q07X3G06MZnZyxXVq8cOs1vyWS
p9X54+HqpVpMugIegSmCXh8wTviUIwaXmAST0qxvl9oeG5GXWQes4rfrL9boXjtXdXVqNh0obhhr
t8W8o0r/wRTeQq3uBQeS4NrDkeOnFss1UF5JJyvgb207/HOWQuyIQAhzsOLi9tOdkyCKAY9Yo9Bs
7/tCs3F4qOV61VjASXeX2XlU1RlkiU6onmWWJiEQxT/YARaCPUygdryZnV1ia89RntRgqEi7PslM
Tzv8AlrqgnPf3dpbQE1lTKt5Xq75J7a0zwzX/HQT8ektBgMacItfVaYGYEklyG1uucMmvW9bY0mz
s8tUqmnbMcsMUKlDrBGdN7FehSouCKhf6dPa2Bq+IdVEdA5m3yaBg0HhzpEVawKkl1yVtFfMyCDp
D8ZPfWAT7iumeIAHYMO4SJNA3uUEl0Nihqn+NlJ7PqIM/WSWbrqu8940Zg9WcOAR5ZPTbhOyQeqO
++oHx6mYf0pM99+Mvg8Hho4k5AODizRXcQwx25pBFf12q1bD7U2KzcCuDCZjwoCNYXqKVpzb66pS
+fPXGBFZQz3VqJca4LCRf97PRrtrs8UwkxDnQGpTwObvmEu177MyH1tBr8pT7r3hm/hG7hQjULvB
zLMLy5iWBDuOpVP5rfFrJ6qhWWKTBdpc980gd0zEPr8dAyAcRPqUImf/iCELpMaOwIIlJBXG0vBT
0s4o+SIpo/HihZrtGnDpnDIn7QHafdo4SoTOwHQPaZgmb1rzD51x8L9IZJNLvttwzEhp+eHnH8qo
mZ75bUdpd3tjs2dMq4+239GiOrQE8iwciW9zM42eDzaxJ0K3MEURsX2wvNZ/nnuh9skfkWl/azGp
aOZVR+9N2Dr7WpnLuNv1+hD0Rxt0Mt11PjUpxWZzLm/ngsNOEP/3yQwYGQyP1zXfdZ0ht7Zl23B7
djxwJkVAwSUkA/uf5Fp3OI+/QlYfmusZTjk92t/sdGwfjHEOl85/5/w81Ir3E0uuErTU71/GcIoB
lzSFWPNKjVw6/iUgV61deglsujN2piZ7i6CzMQTrhSFb0u8oXG2O9gfpmtbiR673Ikr3mbbhLYkH
xjg2AFqFlbRKofZZns6g4g3If/ALH4ixgwkHFAH6hymE5JAxUQwQq35Yehzxvu1P+7RT/iPFMSBe
Psfxw40N2E1G44Q60StKsv2CodQc8v3JvMWvoZKse7Ke4TXxg5ovXxNozauFsBYlIl8vAF+A3eYK
vgO9RflW5Vod2jrVQAefUj3aovSGBkJEXaH5vzH/nM5vwIhHEC1Nus4A/lSreIIuUQiMg2WRXfQ7
w67doXs2vLUVgNV3nN5bUsJ0waXCzuc1husqxzXEUM3kyhXZuhJincPQzmOYbe7vN0jKWGMY8gz1
TtdRmwdMfTT3Cc8j9mUxAxXHwBiKFPc31nkgEj1KDALoXyxQ6GhudbpUdrSoF8QzmLEwsB/iJ1PC
tzabRgScbFnCQsT9J0RRsjO1tcNLFcWCeVqSXQSwUVirnEImji0tFacyMEIuygQSEyvnPaCz0DD9
NVd8yNj+uODZRUn215q8+xassPtMBroAQXzEYBc9xIgGjU9tHDDHLbJ8AR1YE8gvrIKh4XKb2CtP
/2OVFWmBGDHXNUSldEzj6cEh6eeEuAi4JOJiK1ITyRdyc/i+OBFIZwDpz+83XGd+10V+kr/+FwKT
tI4APTwuCpQr6+bxcbicQb5Mo3t+GSlSXV0ENb89ZZXN5Ug43CFScI8GEwJrzrIV1DfN+8d/m/gv
IXEnRcjJBBMtljkQDEgms8q38g/7IOERnFB4Mk0+3W/PkAdsDaBgFuvhVr+xjAeFfE48TxoT9QRL
larg7lRsk2j+MRaEJZKKFuPA7Jh5OkUIJEJ7EIIf7l9GfzumRaH/M9082f9OOxItJYPcZTMcJivA
4LKWibSNa3nXQ1022Tvzr6R8Mb/PpIhUFtUA91zVdjPkJjUiE/NcrvUFQtw1Tyot+SehPddcQbex
9DUi5drowJSHNnhIixL7PTre9qPpdMv0rjmDnmnL1hh+ozWDzO2O+DgOT5aTnQs0pedi7L+nyZiD
By97h4xoecA6D8Aj40G3UCJbdzS+3KA3Luw8Yc1Jjtt+ey9awKtNnJbdoVZrQ/n49y4OPYVvWLbU
CWXPGQLdhs8CJzSRgX4/zn+Dw1YhiAVvZr9WDi7vD0Nz6SM++hHAVWBtZHNhiKOhc60lOsqeNV/k
5mNWvWqzNLVuW8teHXno7/Y0PVgNTN1B81sEJ20Xqs9WOBUvqiYhfCEqVwBEnDVzqQMfuArpnIVe
dyDcp1pFr0K5fbR/0P5/VxZ4EsTzoXYSob7YIhJcmt/sj21rr97Vi6Z0V6PaVG7z2iYkzBOW7KkW
PlVnpYGDch4E2iMSgyBW8KI84q6iSNQAjeXNzZaSG3W8Y1qVXw2Lol6glOZEQinyYpWP+n9MxbfO
Th0HbGpKhq1RCdGzTioqUBksduuzgx9I9zlr64r4wGIP9EhR3UAX7DeLJf9VOYVILDNrJwnrEUx2
W+C8avI5QW6H0ovXIg+z06FHnj75ClGl3Dul5wpltGIiLmuMvbxsWQDTHrZIJiUoZ2tPxqmdy6mQ
RdDi8zXSXvzpvUGCD9KJ1QQ96fXmGAakONHHGFnPA48FsOarHIDAztxbdU4f/yNDPU67qi+Lh5cr
MOgz2PgKxnIlS2uA0mJzWiS3aUwAdnuEigQxkHaY8DBBu7SLJ9UW0pis8dM86drEIQqvq/9d425b
4dhtHGj+zX2JF11XATFJ96gd3tnH5h5eybCcQxfGUeLLXAVF2bme72hfP0sXUsA72rs0QnZVDWHT
PxQXUzOGiR89qAEVCIzwkn4z0yYOmkZCMZ7VdcoTJL4KZSgwQfiyBM3TvNTNyy23+R9SRLNOypOM
T5xrHAXRJSIM0EzjkXcPzgxVEAa3F/ItSy73YbM/bdvAv6XSd/6Zlaov4PkBvah3eDkyPqkoE0/I
Ijirj+YrM4QDKfLjecnV14j9hluFEradYGzu7RWr8CxwoBjjovWWsyWCxjuElUdaj7eDNfsYmTfZ
vD6V/SxFcwLVRgKf6IsllpRzMoZlph7MWl6m4lqRYd9GYqhMkYlxz1kgQbhooxowVQchfSamvo2P
48uzv00E59tv3ecksKHpRw+xCfUuGACxwJAtmWNxQrPJzicFbcoWSbHJsRhKQDqnMblXHtK8uhgD
meP7guLDSur7Dydr50Yk7le5vYPlZ17/mYb1OGxIeLXuF2xbYIbEABHZb3Z6iHYIJiS+bhHaFqNP
VWgA4HHtGnv3+99UElE/ViLR1w24iDPyoch4w33TlHZeLP5j68uqg2z+D+fSuzkk0PBHUGmzsYrp
jrbq6NCMDBXwCJ0lTiTiLZH74GGdnAv8U1WnBBVJj9f2UggFqsjgYkXCw3dafDH4N36IMgOe8LDa
TgVVuEFvJeTxGvqaC4XP7zkobUR15ax6qOk5u4JbdVTrdinH0DpA4pv04NFQzXF712JiymOgzJ0L
H5hdcIavyp7vSH2ugjk6olqOmYThtDB2KCYEP+svyeT/QZrXQDs8gSQG8qug48xbv99MyMKb/FSy
DL8ArxyDxZiKCoKHzf3plDPz4y79iP1+HouIlUwEfmzNvkPZGj6393j1HAFSzEt1JwccGw3V2E4W
UazQ0ka49aHmEg16cDle55HAOxQPN5EKMNovrwhf2ZPE8GydAbCnC0cBQGPg2Z1lM6znwfqNAZOy
VWSyazJAk/s6LSSxFgUj2ZLUZaO01swnAXPTa7vYCU122DmiRKGTFvmSO76/8Bz5PWrLwntRzY4e
gN7savgwAOiXULtF8WO4qY+Euz82Fyestvv1ts4nbOEyk5fY5zWyVSMtFE6OI4uVQ57ZDcSMTJ1h
OBrXmLOYhjR40nh3um8oKXhCf5xxYcuDXfn4S9ToFoq4VOB1ECeimEG56Y8tiaao8pTaURpDBHKg
Yh7yRhxS7m1c3WHmRREqjzsbgK1Z/Prv9qSpbqf/Tl/C2XOHIZsj3RYdH507iOXFs23GoAXZgO9/
bCu2/Fo9u5gRf8MCzATz94QOS46t6pT+YgHt5iJW9iCW7IEtWgwaT+HElwkagVfMMU48f7C0tw1f
tBeqhewFfJui9KSaRDIRwz4KXRKhGoa8DE/tGP7+CTzcgrNNsmnJw3+Ztyp6SKdoJXeuhQYe928Q
C9iYGHlgainN8Hl51PQledCWw2wa+lPpnkjZnmjV8LtxJpKKK7FMzLaUoCvW5in+qMC35MImdXRj
KjHa+nxSC5p+SQXWvqI09ciVsUG4E13lLeI24/lal1nJcWnafAgOBW3GQji8Qf4J8JZUxxmLi/Dz
Pkh5ZbOjW3QP6WGliqK4qcy3Dh1SIexV2roBmVhlkAh+Xpl1y4vb5NZwK0axQJbaexo/cyBQtcuD
MsiJQOUDWz8mzO4f9iRn23U/cvqq8sYIjNh5ND3Ixvz7Bfy7NqNd/voad/en9g44RzeKJd2U1vCC
o/r20KidKcelN8NiaiYFJvyBE8seIez5NhBwqCIIVWs+lV9kCJYkMhMJiFX8e+1hQHwJZEP/bra1
1CHyziBNYTo3fAZQ5UG6koRADvFcR2TCh5AlczAJlPFf90sqnMYPA9WCY1Cj3iCGWUk5216TTZan
101Kj5ap+qOVnNxO6wye/8rR+Chs1PH+VExEJEYmtUGQ0S4/alHmJMoDlxFXMePXioLlZQ7NJEtQ
knxrdwN4eFxWxKjounHgSQxCO9vJ6mZoDL1TT/HiDZPkxgiZ2IFs1XxV7Rxe8qigsLJ0dnDS2xGe
5meRGApYEbjBd2VL+IZ90UUpk0Qh/LU5geZBuZ6h9evEA4ADh4kvCt3k5+5w5Q8uqZfM+xaZzRoD
KRKZTtEPE8Bgae+JQX3eqyD5xfs2muTs6MeYJ1ua8xkZsBG639NAuAacTSYPFYb0fxmmtz7SzJBP
1gHMakDg4pA4rsTjmBQmCQQmVAS1FV41wuNawWUh20KwMnekAdapLO8OQ7wLtccLbb1YoG48iTML
iR4Egcfgg/y4ofDrjErHUfttNPgG9mtyvUKm7WI3gXt4QT9E5hZ4SimoJvgAJS/fUjCnEt+ysCom
svmM+kbTYixPVSxmQ/pEI5nc2M2hzRQR4SKdMYTXLNSW1SQtKuV4krR40CaVrMtK0/x8OW5xjINM
MaZ7nILpWLAOVbOFQw1u23gFFzFdg2sk0CiMldI51WSAtw/0cWQn292vkoVjG5Jhwl7Umt8hlE0U
W96YByaEeHc+mjb3Ev492uRnXLe6VhwmLw5msTQ6hSeIat/7Ru+BqKUto47KVa1qMHhf6ljTi4pS
8OlAFc2OWhsuRIsmqrwaw5tZHtXPqlQeHuBGEFko5tkYzhhQJoJlJcUV4bBQ16SfzFUnBDGiDWY1
DdVuUcuiCJOyiFv+tNDdJSzPoo5p/6KKUakQp9ubJeIDt9FKzkC6JwZNpvUojk0zDmXOIHxLz/TK
ewZBmLRHDKFQaaSbCi3SkUcWxP1s/EqbeipkqlSN0f/nHadKHT2ZRjiPkX+HH4DqeUhbnvSNd4K9
5jt7mUNUjhf6rX2P999/RaklHh4hQUofeQDgQ2elCmkQ7hXEjWL5z++q4f3PyTfCnenCI2q/61HZ
87TB9xPEKAk2qWnaYomArz+AKcgYKxTQyiY4CPn2Llf+9TdQhxqNMuucJRVj8hbg+S4s9CxJGRe5
+EBy2ZksYLGj2MdCE8FvVjRJfyzfp9iUQdf/Za3uUZz74BCcf2Dr9UlAn+Q7GlhN3fwsZUPTUExX
B/Q6bb3abMIaYZ/JRgOUH01Np0dkip50r+6N4klcCwLw9NUGV0QNO60pMZHt11C9Irx/4iVzAnpR
k3/ZpFQvxWFLCUQnbq7LJgXRiveh3L1gDoEBF9rsbJEB4t1/C1EaM5p69mChW0DYDlmAiDkU3cyw
HkM3kMNpRBvp+3uRhhLfyVBUeegKpRTpt7IjPdkzx66kE1i6hZmyxSr9RjuhhTueB2qk2isx5rFP
Du0xZ495hTmpmGMoytWl7qibYmEJejWx+GLUPX5B3oYC5E7lpd4E77NaZiJXc+njFoL2kTJ9EAGn
U50cCgdm7V3Q+jRVC65OYEc+emsk2hY9x+zFAjfKQH8oxtbGJ97DYA9+pB1fxfj1BpQJcWvCkxRf
6sPYpJuX6zN2eU+ZUL2G/DTzARP2kAjn+t6tEQESGjlCeGLsVwc5R1fiHgkJwPhFXHfIiTExcluz
zg6Dzs4lxJK7ieqVdVRvbkRRp1Avs0wWm4pwkDUSUtwRcIBsCzQ8lf+DEQ7X/3aeP3oPWe5oyL9D
RGgjQaMeQA9OCAuOw1SY887b+Ev3VIoJ/VP53lbzQec/xkRkzpItnZ2CeNBYmcqceGe6hsnBiKFR
TvT29JL5zSv8fe+HV/+mTdudRb1MJVEi+keK3OyGGGpTkgoIPfsvqaUfZ2gC2pW+47tHwK1GBusy
yGuSxLaRo8d98w6djE4OLdFgadk2fKwqiRNVmJrgmSBKHeQpjmwiV+ahL9fpgrXKoJnONZExgFhT
k/DLgTDHGGDJOThcmbkbvBzxSizkOMqiwSPYsVFR2wreP3FNPOHjIPTqNPOJft8jInZW77Njb6hZ
Ggu6S6jdLpC5MrTMdfnZdLHGs/C8K7vsKIo8Fkq9GrYdh0f4suqUyJ/AFZqGcmFQOGwdoDxSH9pd
QNJ/w1Mkkhj3rFkKhEvc5V1Hl7oAri5MBzsgyDV3OA1WmDYQUTT4vUV/rIe90d5twk+4jvBn5lPy
P+TH2RVAl8i1mnHz4uohaJ8R60Sk3a1pL1DC6EFvptHSxzGMXhcH8+iUWmXSVkdFLrRiuJzQMQMw
4iqTiBeFEOPrxpb/fgEnYW7YU6g8KkxCBcz0/YO4dM/vXAipHWOK2jT/lJ3vay3FLR43awYCouWK
wSNhUVu0jyvxNF/XQmT50rSNEmvB0jY4NhSuFDdG7GfgIQjiZHVzlyiTqaYzXwq7B4HT564a0hsX
06aoorCAaVK4fy41imEVS1Y/wLUOc6/cHoi+P5ec/M7j/usn3nc/9p/mahZLVyQCKE9eFi5BMAUK
aRVag3NplnMwTP+mvAXCPx948X7wuWrpKppXOiW8t845iwkRrzUH1uHjX5myqnCUudJ35s85zB+N
pBHytSgpDfhjXyYlSXLhh6Z51Q9G/KE+N+0Bs94Gdmg8b9Zd4Ytzifhrb5VPYKabmZnYQq7NY2vQ
u5Uw+oPIvdTDfu0dm0ctAfUJmJ5438Pj7YC9rHVOTiujygPMgrWqpMeXU0uULAqB4uejlr4w9+eA
tRH1lO1tvMr4KGkVxwcDcpu+EA3dqA8fTW40Q79KPQ+JejfUx98ELp19Cpe8pDZA7//kxkFT7Hyz
7vy36NMWONFaw4HSzDC6EDLo+pD87OAKQQg9aM/ltpOshRj7v7MxQmhiZ/jHxg6ZwWA1CBRM0imz
18dkQEulVeg3O2260V9g8ww1JiqGXaubDSQz007U0eOKsYkNERKhiDa64idMwjFu/URQ2gyJnB7+
0YmcjTO5O3bkRATiaDQcx3aVMhxvNtZjqoUC2JAQi2+WlVezrhpXhp/mccSfwL+bdURds4H7ht8O
yo91E50EJw9UoO1qJR7YGOw42IoRXdZi0a9rayhuYgzsTz/RaynXUmF9aXbEXbwmfyXsbDyDMe8m
vQmMsl+D+5qlM4n9YbWCjlFWNw092WZ3RnxA3gCQKgI+Cm+GY8jZyX2o8q0+TVZyZ31LArIdBBUS
OCtFUP3omKrYhIzs8P56gvILkxkx3IZgD5JzGnog03U8yynmRqBJ2uZlbbyuNf+bKIR3OHWmH+kW
3XF70J2g/zoXSIL5eOe/U7s75z/omu8wzGjZGeBaTBJRtFh1RVc+rEXuCN9bYX57EJzFim++k/x7
VVOtBxPov0GsErxoCVBca5c48p88+zEKHuU0oXBWJcg7qwUD7oOZqM0v3USdnDdpJcBRXipajur4
Xq1hm23Evpd9bRDBbQ5E9r7dcELJF57qAQjx6ziTeuJytmNAH63bfGvcJ2aJHgWzWXr2cwvhm2uD
IO4g020BsT7VAsN6bGypajM7QMppIiLdcn044xW8DfJ3AwM9/1KYwc/LH4Kc6Ku+agOtGLj8tVq/
+9b86JvKfW9o8JkxkZyv1kXla6xOt1+Hd6WRUwv42qOMgRadzJP1fxqdVujPW/ZkjZSHTsHAD93w
uOl819j+A7Tuyyt11BVnnPq0iLSxb//9PtIY8pGiL9ERsXfOo9MrQl3NzVNFsQC1GvIJh7CqmasZ
nvt++SwMApy/ZCjwl9vG8OqEFiuHg7jRJKpbtaMPXgCOzCLXKIaRwoWq9pC6PpneVS2DzSlVOzbl
UGpTYM3PvyIAHfB1uzqRT/LMNn45Gd8Pd7Bs6tRXgchVdIjx9gTLDTUMGceceR4nKZ1dpbCIh5EV
/sVD+waIeE4hZOQCmYUCR/rbaKvfE6xzi3o7sl7nTHPRb6j2V3/CJLUapGvD8311/a9dor2wCWKP
253zyNtgOJnoTD0UtLeZbg7k3LgVqq9wXrr6K3U3ig/yiT2ga2pzG/9orq12aUYsjMe2upxeSVCx
YX4MbvLInhbSDi2UCk6bVskVq4aKn/8PXSkfOCbjzJYeo+mSbqeL5acTWtKmByRnxdRnn8hNE1oI
jZNXYKGEmvCf2ZSlCf/yiSINH/8b51xdHa+hEgVliHJt2/7Se1TB4l4vGj49sGvsD4D38InaaK4O
S5gpCWzLX6wo/YNKrpBLTP3ZTeKolVB0Dz4fxHjEW8lpN4mbssWsKFgLMjm5VhSWAa2+m6I11+NV
YFgRuKxiAX1PcUlWYWtD6hhqVLfY5AqQRJ67OpteYDioHwn2sX8FirnxkqgYU0d3u70GgZciaY9C
0uakshfGJ78hDnaqWifm/ziRtH69Au+uIKkILlVRCsvuxJNv+0K656wEqmmpgAfsR1bXEWysvjBy
JlNG403FMk1s2YX18itzocepTrw4Fqv5TS2wUhT45V6oHzYhoQ/8RYTEFZk948Ao9fgY14ftFwbQ
Ph2E1u9m1GbtmvV3GXoImN6/7NtH7tNy5qFddm/V+nymowz/KrsuC+UlHXKkffZP16e11ouBGVKx
80h0zJQV+v4QmAgbqY2cwcvWwB39VaLvjkBLvKiMfuZV7CgONpKhtYwedWZc8oWEDvvRAqJUD/QT
FUi0lKU5Oe2HaxPfS5vqfyUvQsSN3zAaN88s7t4PcBe5/6OB20u9KIXsseAjS5wmr570Tjj+JnB5
9K/z2jPW8Wch46x6Zo1U+R8KbiW41B6am2rbfYCk6Rk5Z4V3xVEGLsA9LxnzE6XJlJIFPujhraL5
lw9YJDtxMOah+rjFda9MhtsW3VGDFS7eojlhc+ptj8qngTBLkzWQYJ6bcA7tlPilZYCF5JuunInW
UHm2VZXp16Qfoi6Xf4XBFla4CXCkADJ/WlNabOoE8oqSKWxP4mNTbB6hFtnE7tk70TNTSLg3UZtr
HLw/+vFzosOWO9RIjPi/Lj6D5pkrQMrMKvPqozoxHbU5e29S7SckONNQHxCWosMnvm6Pp4YldtZe
lBRG30Q1mJj7hwCrMn22/rSaQE+mZA5P1vomaZ17oelGtV2QZdJO1wzDOfQynI7Nxon9LGmElHZd
M29GhRc4RufuPx4o/sn2/XlJL3q6B5DVTauQYPexv2Drl5YnEa2AiaeUyOXUnGah5RpEB5DKgnzt
ufYT1UckzcFBBowMhaZj5Btc4wvTc5Ivb7qyUZmPC+tIO7Z/52xOeMCQipjIxL9YaQxec1tXLcpK
T0V5rGjpRZIFqWI0Z6tnekeYDMpUueilUdUsQaHHq3aepOEIc/FQVcp63IYNv2x5QBmx5D/KrTVP
zjXypA4VR9zNlRQAD8+Nr/MQZVzgjdAxmg9VZyGmQHo19IHFvtXtwdLopHVzdOPmgFBaI5RCT8lT
9MJJY0OyeOnCsg0swSg3TcYLI6maoCZc85H32ceLr/ijn/gdfRc3uAHm3kAOeKtsc16nHtEmkKwP
ozR8TUbu3/vzuNqsz+U2snI6soE+t9kT8AUUBcszfIOrhnSB9CMpm0uRFKfdc21suUoIVpBp6rEL
x2xUXenSzZLj8znNBOkb6ay0wjgJ6jiRBA+lFJqoVRFQKfEmbH6K97Ie2f9c4Mg7nJXVTkMzDmFH
iZDP24plJAIeSgDX5D0uJ5x+Afhj00OPxGrbr1x/7Dp1gVr19KSOuxXdxgzTGxwoUXWYwofcvMLO
VBc4TM50+L0UYV031ZpOvTpY2Mj+BQ89TdxheEul9PV+3Oe62I4KET0vH1CCpS22Mh5Yd67J5qQ3
8UrZQAN4vfP97P/AwQIpVyfmN7o9qTHaqra1UDVgQeEividxvVkvskx5v3HkQ4NuzhcMce66gXs6
+RMTE5VYr2DFPIc/eB6l9yrX5p8bId1oA55Uayl8oh2V7roo8SU7tuDYEmvleNUKIfkfdZDLUx7M
HpU/mC8G0GyccJAMuM3UV0GJmByn3AYV6dg9gOZhbOfPgZRoFiWaUXBNafPEE16tkE7ed+izfJJz
IbAkmTM6Zsz3v93RQDkhpt63V5Hz5mYp6WL+dC5Q/Kb+Fq26VTuFi7xVAvB6YWE+87MgcmDEAve8
Wq3BgDMSnKXMAE5v7ydN9065RSwLtz65gQeDfJrf5pwR7xxQYLOK9jUxY0Phwh1R1twGtjM9do+4
NDwNUZDeOJqwLTSmHcVwWo4QuGO+DyZwdODD9NxRSnFfxYU5zCqnMVa4Pr/emwb46/bxPeVHVasj
WmwfatviLmJ/R6pNDMmsQUrcs1+hA0/+CpxR7LOFzuYKeaEsnasIMXfwqD4l+baO8Lm1Fttfis4L
TT/PxLZSwxmlXRV/vIWwAmaIGdbP5KTJqkGyRP2k/is93q5XpcZS2mMKVvjxU9saVJwCkxYAoxOY
/UBSHRdZoqnSIruGFngU7HCuIZtUPr9zcjt+pcIFzvySBcLC8rUd8nPOF/DCxAfYJVAW+ru5TFWy
VIYsfDSEc9A40OQMgBCSSxaY79VN9gHyeTOcJtFVdDcSqLlNBl5EQjV5OD1YQs2/2rOducMlh4xE
YiDBZkRzQGF6M8IAQAKxRNyjFCWHjyQDmqJSPDrJ6sjn2FU7ABNSfcceTrvwJ0MY9EJ2Np7xN684
eWtsskYB4gk19svOU56nhuY5qO/RJ0WvCVcu4w5X467BFmYZVxhypfBZniavXHrV32e8PuEMRTpe
7v3oIrpVec9WMXTcoQRMnn5cs4bvQDGAIoK0DkGEkw5lkQhjOBPEQSBvttqGlrwiWHAzIp7X2HHp
I8eTkNoOJqsdNqFcapN7aK2EPjIKEqq5twI5HdTY/dyAGOwz74OBByPmulqU8Q3tzHj4NetY0cUr
NahMDrZk83VvLvIlYmLBh4cRY50flVK2ifU/n6Lnr5C0rPr/4G8mx8DV8SHORRt+RtMdyrnyo7ZD
jAkD36NVz5EfgRwMAEZ2rTQb1HmrjQki9VhuOOPLU+8Ldhkd0dJWI/9+mPKhU0rpgutQ2VhUNzYM
VZNSvJOqkydSvdnnI4k7d1PxksofkyMmFMKTFkCDOk82wpr2bo2D2L41RgMNCooVo5GqUCBdmAEd
eOqwUnSTeTM75/3skPTMdW1Fp03lWNE2ar+swFB/IhuLPjSP1AEnr2on0OZDDiXo+TDXAt2c9EHV
ktjkuo3U8Nq/UCf4g6M7xvmOJHkIl/yEXwFHqVdxG2BdQL+ffuZlwVRgaBMgDq/nd8deoXhvc9c5
dwUjH+5U61JdBGiUOFsRSbaGsEZ8HpO+Gm2qpJn/iVIag/dGwoatxlrbSyjxTl7aDo0RsWFTo8c3
E9hlPSORD2wYW98Jn4k1Wn9+iNcg3W8oB1o99glTNCzIX5YS+YHCrr7+mmkIiFlStyGdZeRaT/nd
8KD9zKXrr0OIPZmN3Dr2ucxJaRcHNkA6tGZbrVOvmYV5ZcneIkmwjaTHULatE6hBwhSBLf9rqfd0
KHCHBDq62P2rcyMhEdtJHE55eqPXns12SqYQEzPqAcDGPTrjlvRA6Pv/Uv6KPXnQL34xHL1cjaTB
xdSAp/7I9sDcoVUB0WmIVmr5JRPoLuAUzQmc9/krzzJ59A+Hh5jeluSu4i8LDSIMya/UOznaYRV/
LIn0E1S048kAn0lTGR6Fle2+3C5UHDVl12y18A4ex2yrcQzj/u6ZGh6SiqRAMWY/HVFhUB1SLm+5
ARHjUxSKZtLylz8J/UKR6GSzgHCRL/y75Z4Bpo77W1b+7gf+I56c5TbDkkV3CYM0cxn74ubQKF9s
teaq61MZsukB9DjCITDQPTgNp8KTnpbKWE+ayGg8UvuTXARb2LqWcsIOy+3izgO1ZBMvs1yHm6//
Tl9cza7cBpuLhF5MD/MLMy5JmmGKYKdmM7ivhPVTs6vVbHncnLjeL0+TYv4KPo2IaWAb/Al9u316
L4JuivT6XZJc5/fB0OLGdDJrvLmnFK8EJhwBqvC4hEH7VmoRclwBFYpnW7KjCh4qYIKrJjcQhz+N
YWx1DjrfaSfI/S6ZkXSBlnOVoIMTHAHJqG2C+ZMz67DuarJcITJf3DawRl/iok2VviSF97v0UUOm
C7kmH5CDXo/CtgNXBFRz4QVocgv7/9orL8oKSx0YqBe88jspXp2wEFUU/cRJ49KVjPSbCZzPIOqc
1FJwB9eLrHOhZJ3CKmeJTsHsvgS1L2TbhfsCWhvUbyQubYNu2yGelCxLRBuSF2Vy+6SNLIvLPw4W
YyzJsmAyzh/RTWSOaEefZjzsSN7mXvmHcbB781WC9/5nn60AlvIEGngez9LZWMlZ7fZiK+INQy+h
Dav7NyuMHicrUXQ+OEqADesOUFZFVCqSYduJILWESn2Max+wTiAZnz18CRQ0uulpMydD0/ztEQ5Z
sr0Lzs7l84ZgNIUCzlt2cXbGd36FVxwNfSEct1cwlphYaSqzMP9WC0VNmNXREld//YoGIPl0QxAd
Cb4Xjq6AymB0l8G3TvZreSGryKzJeLnTxbz46hs9m02H5AFniy6rTnoc7QvxHg4ojkn9SQcpqHNp
c7Yu0ssS/04lDJvEWaYqwR/Z6nFAn9uMqTdbIhp7ZFmM9MYajaXQm7Vjp+IAZzdXrvg+aC6aE7gE
itnZDdekyoWkN65gVyAwsQd9Sr0r5hwMQtZ8xZfi0/6fzbaAr/XJQd5sGDsrgS9wSm6KMO7Vy1kw
AbQ2P9aWOTtkuy8ofg47YC/G+y+m68aYSQqDmYGBJ2B+811Zp3dzxRB7Aje9ejNUhu4Y2kKe+Y34
LAhdOLCPz7c/tbKdoZUcjVDLYrHeM/p8/XWqF4voZuJyA3v85SvSZSOXursQJlYZSdbSST1hMj2W
g1bSBPqExzS6Vg5UQAIrjkRnRYDp7ia/ykYQrM2Pp5MYibtSdY+VfqIFKkGYbeVP0H6iPjKonG+U
dAfemJA8bAeYYctR8x8mpkc3ssod1cWRWLsHKDX85lG3GZFRjQ3zzB5/ysiPXpbq3mmt4kuT3Sf1
9JVngG/17W1z+C0U24POAwKSlWYNio8iNjC9PENYmbKQene/g1qC9IejPxXSu+wCfEEgZ4Rqmrmh
/mOk+uLZpzkNXryJ1X4El36USZWaRkRvYTTstXJi40ntkJChl1wxRMS+h0iuE+XRJesP2sw96BjW
3E98rUT+pt97VPf9e7SPULCbLnjm4j6Z30NXRiyrSdB7dX3f6SVonXkW598b2nGs6urqB0j93zG6
DD4kAakpuFhrzUqmwVngUvNVhi8elNRS0uuQlOqcCcx4RcqXML0nHXyEdfU1tUILL8GD/LJlfBmU
BOO5vAaNCK0fWyEBGkj7Bxf509y/fPGnusD8F42L/bI95lBFWYDc4CShuYsneUVRymcrJmOJ0jey
sAaKnErM07+LeD2owFMvfhzxsIAEXt//maKYzpTGqt60pJMQsL7SNYN8DXRtuAY+clAhjNw/wYiW
o/QroSg6to/8qsaWsuUzL0n3CSd66o/ZatmDdF9i7a3XA2v+Nmr+CJ/VGan4U9V+ExTSXp1cs8YE
ri1vgpckN0aYSzT3KfnnsguEzZj6gjWb3HVRSfAnxdn6u3vUaiiZ1ElM6kRyu0S73T/hYYrp1uOp
2zNL+CEHHa0f6WKZUqiVOdWfbFkh8pYoJnXxeGig8wQiDOXIqxikwVbWxA/f2HiXLYUjsmhvDueY
rU1Vm8nAwuuKs7K4BwBcU8cOT2BUt9HjQySurPMTFlwz1G4iG/pUJFA7eAO1Z0rle0MI7sWuQkUC
WO1T+xmxA/jTdKPDGb43M5JiGAdH9JIZZv30MzDIDhiztWsD091Fk/q4eX/CUJRKYCeZmbcFUbnT
ff8vVYUmSI9L0mP4SVcBFhBGcQYJT8KjGnoriqkzuOg4cGWgcaOcu9khgqAY2NjR6x+FWmqAUHVK
xvP7zgQ6kVV4QUKwhS5+MkgJDFt9DvmUuMRslmOnuaKpr0701gZtAe4xaMy2W2FvemfKF3KvjC4A
Kv6m3WkM5YgT+8Fmsr3Ef0upzw4HlBhvpoiuqGn5TfSvHfbCS437VUMlKKqaTOuFBHfDxvzO/XVr
KLlYHs0oUjhAMOgAfMzYZtjgPLLhg7VVxsO7J7pShdxy8sBvWzxY4129JJ1sYKqaJO7dSVk8K5Bx
VhVOwWk/pm9RkLHtuPbh3HkcwwoAXzHYinebk7MrPSAy7UoK9HIxwwOBScRQoE7p+UNOWEKuCUqW
RgakSkGoiVVRIshC1OO6sS5iQKJejxHfWEP1Q1DMEFos3mc1uyLQ2vx+WaaCWZB3gKKn2rs5hQq4
LDH7gF04c+YHCsMlAYogdwvWdvuYsKVa65KT3QAnLhX6EbYkjzAqxpCX6Guzk5ByjhBcb7FhLB3b
F8ADPgjWZTHJlJM4Tj3KEgGYY5KwSMTi7PhUhHpQ/OP7LY4gymfO4xRWuVZGBvYarkC525eBsbL2
KR7hQXjeuq8UzimvPJlxq4HL0uCUKUZ+jYAFFIsRYcK7rGHWIdQ6OWgaW4HAtAbcwibn1u7TYutd
rGiVmQ7G9S74x7akAOxqlts6RbZzQPHGOo8MzLDa2t5zq9mXZqILEhHyX4rcTXKMYQAHq3CwOsX5
00ebPMq+ZrOcqTeaXKxEazTVI/QRrQpQuIwkkOjAqtiu7oBgKqZpBG0nqXTMsTlRkB+lnRXthGO8
L5cE8c6Fo7ZFxluSYVCidn/Jftail7l8mDe+NwX70f8Sv/oHVbvzwxXJADK2mtgS4g+wvCD9XZ8k
/mmuiW0uynnd06VFS3LqodZDDfWls5wny4MnWdx7cacQdXgxIm6ekLAnpsIBkBWfomfWYcH4FJdj
ihdTHLG5NvwGNgsYlx1Ww6Yf9f0TyoM41v2Pqv6uzHXowov5bmeS+oHPwMAh3fsTvTRmVXqZ4mS0
JKwPGQb4ZFsI120vLAWhG+7URWEjLliVtS4ewfb2ZNZngWC4qvzSrZ01Czt3tYzFvclC80lWqis9
Q6xYW6jdP7uo/3HKE2zQIi7RIcIU1WUtAhj5f2QsrChy/iZza5g6BdsI/EO08U44/XVrFwcmavU0
bfT5YgwWdLS1QFV2MO5fAhd7C+3PGsPA64yXuvDAYdlBlrRXnMv9kZw3nQb3B0OK+iOLRPCawILk
LmzAGHpkVHA/LWADrpw3z2cCMKp5V1vlM8OH12p9XgDVq9I7sxijus8ni6jkW5RggHhOJci/iPWj
qEDIgoPwNsWrpWtedmbba2R3WgUiUdT3xmUaqy2Sl5x84Pylm+TZPmEDqq52Q2+K2vsALikxGmlb
SDFhjAz/bebG8HpRo1s7QR7ohNI6XO+9VgGcQamaHXAHF9k+5kRAEUNjolcjafUKCcrM5h6wG/le
lxUdiYupy1eeyip0L/i1xFoSo36ZcMy38/CGlrybbGugpG3wHEZiTjuXLnofVaLSZJ+Ye2JG0tjC
YhT2UgC69eZwzMYW52uC2q2PtxjUHpIepZzxPNY9SvCSX/sghDhcg+6gsnvNeSIX74rXOtCIj59y
6ko5iVb/Pa/xfOwdcvffAHlOzL+34p3vIk6PvE4EivBRTR9H4LXFB+psZZNduqEZZ7FD2PePQu4D
9dYP6MksdYavxjVuZBcGLpUkI+b/cv1gH1C2Wee2ZvDGPkpb+XFfRr4Mte25H8hjBBm0H9KIWU3b
ON3vA4B4AGiWP9I/V/nuXD6oHj+hCan1q/FnK2Ee1ObYDUmzqiogQfcPI2U4PAkZOvgz6Kw9lf7o
46db0f8g9NofGE2z+9riopphx5jPokMrzmWdXXxSerwXB1e4poj3fGh+qyk910ERlhuBGWeikrsb
GuhNbSW9Wx8og62FNe2YMP9uwXP9ZVyjn5xCcKXHUJtESnSl2QZd5uFSgp9WRKcv/x7rTkGnBi/a
VUkklbwK/QYp8Zx72jZNREuYjo9RUjezakKBSvm+BtHVHINEDi6sP4pw6cED0dcAZiN469yXAZ2d
QCABqWVDXS6U+GbGwhhnn/jrvigcD3pvx2GCqymYAfAi6fBMe5GoKGFxU9ByKbDbqiPE5ssWY2P/
q8b3OMGqt7Ym9EsD720eHbrYVWQu53s6N/EPtNrFrIA/9vTTbYp5uMgILrE0U0A++TVMZ+A09qWD
aHxXWqY7y1JP1oudpdcQUK/rx3jBdILnD3E/v1pRHcm7MiRP/eSwwiTMP8JPlVkqbXuYrgaK03AL
fPyW/Y8Snboy9uE45X3z/vCtEtc5gYn4CvA1r9ddONvvqiPe1ky/yOhpnuKQBRLBUNSmpW4LgpV4
qu7mGeFLkWfQn7ISbIjyl8MEKwh40a7yP4+dEjYebLQzLKCtUKRPbuZUVlSdCOw+2E9fj0yA0euS
WxBaSumVcUt3Hw3GzzdItNiVl+lcFH1NTGb17oJgcVcZfFpBVToKEAAVhkT+FT5cWOuhdqnNhyoG
HAoQVmsaJhKyCbNF23Bh0b77nRDnJ3f0qFcUe6Iekz6GFbmT13CBywEYxnkI5YBV1WV3CjpL5hmh
Niz4FuqgG3UKXckCujx/CbTIDFm7tUGdbTOEaC+QtBItuY9LraWYbUvM2MOLEjs57zGgqI6snhQg
en5Qlu7HUI7RHRpPj6ogAmXm/4J33VFt5mjQk59Xg1onWQ7NGunWWJfxsuSRotGImIctk/+SChxO
sWwFlDD8dkU/so1jommb9ud749kojX60AflBM3DFg33LGMrBuLo6w8D5FjOO/adFJXknRRLUey17
N4ZJpfYQmLpZ0CS6Uy+8f6qgQYU/3HDsHWZ1d53lSbhDEnBHn+fyTU8/4/OSsD3WiPtsO8SyWsfd
QE6v840vMpP3UDbeM/gQ8e5JLPBv6XnpAvE3YJuU6qXBjRg/S+siR1OBnPgstD095jlUiHcdmg8z
Yb01h5vNlDwxkB0JprQWUBusVnn4Yd0ONbi9G+kwwz/hJzfM2g/q9p7zlyZuO47aUplqkGjYjNf/
8YN5F5T+DcFHTuE9LJX8ARx3ekdbvi65v/h3kbS+1SFFnh3MCKsZWdnYEOufu137CzUOqdiZ1H8U
AG2DjqeErAOqD25M7rKzIo3AIdqpfkgtkMFazdBAwzkf0vCOEAt4qY7+7aRIHkOtkqbDSmbpTYrp
SLKR9uPwU5sACNHqiwsXlDVrFbkifgKJ1wq6cSgVrvEqU8+B0c59AEaInvpSgD7iHt0SqwY5EJ9+
YLXUiOpPu5n+06HqvJvGxr2OH+LUhzVtZDiBOSta/hdNamTDPtQDeZJBZWde0WqiBh7pp8fJAonA
X+U0NMBEnGeSR0sTbvJuXB7LNHNpiayg+cNRpLV7eIw9+ZDgSL90NzAilswqVeYow3rkMIq7dUca
8iBFFOeo0xJ9N7mN9pPNxEh7GrBH+YC6fkbl1UPWRGoFLpRGP/MNlZjbZhHiLNlFS/gl7t5zEdMG
7huMpqbkiyI6nOO8H/giGsUYux071zx7/nQHOXW8UoN7uum7iMEdMvtQr8hnq+kKqGGkjyfeek6K
HWnlROtxRpXgAF++A6djqkRjA9grhFBFuDSqEZt68IY3e5farL0GWDMXNK6pY6cUzK0rsqKM2Xji
cdn615Ain8u8eRqa3oSL8x29+6W9y2uwUDbSRkppuWj6WW36ra/bir324Y44deo4+e8nfW0unGEg
VJyN4JgupszY6yMizruCV3j4IdoaC9OUV6qTzXsJXIvOLqhN1XYGtFXnBeUx8LprOLtN9Y9kwkzu
3cmLSIsq79U5cxquNFA7MpfFE7xMOBsaL2bF4DtxSYOg5BHqLoMZYlfs1Xx6rHXg1HnBQs1yh2Hb
sLxKeFbZCjyCggEqRmS2K8nDeou7pgYASunb+kbzuo32LkDLzYoXnFxH4nBayknQuXoYJTpxlOT4
/TD9nMcKXrPkwI9mCsOW5s6SBdjH1xlEAysxpJrgXN6tpM0NfLW8a6lWDIl+rDzljaqrUv+q+lIP
DJCVtApxQujG5dS6sol3NTq3BjgR+XsOSCy2xDU9mcvlnDY4AT2KZJ0hUtfEbDUFidbTXtkyv2Fl
e24Rr96/OHM2dbhZ+2Q86Lb8nYEQojNs9epiYX1/F/NxLvtS+s7fH0e22hC0NEZm55EVHIFoaHue
/c7Xb0LnjjUICo2WM+KmzZSSiwGjVB8pnCTD9Jhp2csnxh1vundd9BgOLVOYNjMqwty0KBZNx6lf
FEbMXYf74Y8EPn5VcEqfHQX0KFW518wPM3pD51TuYDEWO4CMcBWGsh7/hQ6/8MiVgQVdJe1+aayJ
Ca6lcqlN7GNbPKwVU1ENq+kg4p3DkzN/9SUh86iHa0qVYCrumcj5hPX1pCZ7/9l38r4V/zbUUp+H
wAENc2qK+3XtFeud13zA9N2dhN0QcSVeG6Q4+MyhGkpk5AvbTJCrS+GTpkGLsg4zbzD8erMBX5DV
J7+oOKXMUgTjNFerYsowXiyYw1z83fVFrFF8PsLKPGpZb2vzvmZQ/jXq2bnVzwwHf582HUmDc4qV
KE8dDHGuOvLrjndtCA9Kd8kAdAePKk0Ez5L1BoJj89WtwpEZc2CentxbU33QEK7Rz0jUMurcYda1
hN9KMlLH9PNWoPvoObbu0p1uRnBS9oGZT6de3Mxk8P6oXnFnX9l9VcHrwH14/5P4KliMD1EqKPJF
50W53JlsgmNsyBmFeJujHIGvdbTNfHnD1KtIO9dZOUQ11fcmbSPaKRRvMpZNduMc6AKhxua2BVxf
g8lgffFqFGvq44xZ8UNWNCBWIzlV/KWY63vj8X4ocNSGc4+4dWp7PFCFzt4S3a5pxckNlHpLvDBS
l+nqOGBn9zMzSAEjQ89LWBnxB0YLuf2wwgNbMqCBpgjnpNs+4iZdpwCNfJ598CocOreAe54D5TSS
EEWj89w/XThX+Bv2I+iGDXjRD6jxH5duG4a5whuK553zm1dJk4Q/zsH19HrtgxT8qQiD6SQ51dUk
ZQBK0QkFtVkLMLQRfLYGh+bOTDiCWmtkdKEedXLOZO/9LtPeVJq/bHIRUjfe4V4oJqoeKap0xktQ
DIMbCvFIZVOI9b7GnpmoVmKo+FOG2p9T6LyGFN98sLo4wVoXYXadpS1VxSOUraYADVAxp2gqotoY
R69cH6DvMkPdvNNzDOhvlcvloYCUdlC/3FtB46EnaK+bD9ZE639YsxLbpONopReLbExE2RSQMX1q
EaddMQeW3cTCnF9QMlOuvNc43IaUg1zCsfgaIRLNeZ2nTXF6V7hClMpT81od/YornUG6P/pE57fZ
MdJyX8UVbHVgcRS+mEWVP8ZYGRsFqg5P2p7i96euR6cBAnM0X3Loz9PaC9HdVBjeQyr2/3aBtKoM
szyG/NAH589Rhb5brIp6/9Isr67tISxInekSixLPXnBrQ4izUIdFdPx1oPc6RFDYK2F5GT7yVlB6
LQQUDC9jqEiTX3eo4pm5KM24zFzYMiu5ygrJI8PXTTMNJHyOcLY9rv1c4jSEjH7TAkXM83ySWhlT
CZ8MWTihCJqaB8gLvjz29U4wq0cuoJrC/as5+/sz69GevjAXdxDYvXAK1ucvsTSoSvJXCte4RwaZ
YKYNANCwWi5m5VCt4ZPPaeN9SjarMyNElGN/ip0s3Q7pgxMZXdwdcQPp2fiQD97rZuujg3kIa11G
CWxDcXnp0Hgk22Wx5UDIS4/5Od3g2ogyPeOoErYKLXFK+lesUz5pi7tN6/l8U6FnGAwRSScti6OG
Lg59FevCpvS7QMp+/RVtM8+EhwIFWjjpiW5VPHZQm3qQCg+amYARiFQYZghVkQYwJ25cgnPsykRu
GKVtDMRbLxkWuaIUccibs1kP7MW8qasdc6NKPTl3e26BLiNkxeYtQZCoCDMSFHo8k7dzAKAUH0pf
86+JT2dKlgTtK6Ryn9vpOfh3QgOQ1WjYEwqRMiiPpX573CidY0tlB+SPCAl1KrLFNF9eyiXxE3JB
9UA4nZPlv7F/AZ3muo1VABC+L6p5JbMuF6jyzf+4ayadzbHM6+cPu4dAb6x1EBseCwOGv4zDKjHP
g6hryBA4CyfISZ1zCqCFvWJCT/e3sMCr0G/yYmy5RCIwmWDITenUyzy493uSY+NZc6lXH2R+8Wou
ZGGQZx/ITaQOO1TimH9zThT0Wf2IUy1v9pxWd+d8VG2rZzRWBl8dGhyh4WWl5cO9nM0LbWVALFvk
ZDIpWBn/eDtKyMGCwdjq96m8B7RG8Nuo4CcGWE0cTlQximdkXjc7ONUAvyb9ADJ7G8n9XZYL9hVl
8ZMqxvaU1LzFljcyCfvnUp0y2UxE5IYmT444S21D9z52K+C9Bjlo7eXuAj8s8ctkFsOFNYgJp77a
eUvNijKM3OhW9TjPzayFwBu6zxE0KMoLQXCHOrhhyuZaUNXbjIAK/5SJuTOplB9mNUmXzedKlDp5
/AkNJDldpYy5s3VwYm/kpqPntI4qbFQpan+mr6pyuBuGCIaQdFUCpkVWVSTt9ovcIAkmbkw40a4n
5m/vvhnmKanjk3zAAH3ejxP9mst1XwCwDXueMSFGWJuwesSy1hyC/tU+aFnbRHBAEkxRHR/U6+k7
+1g6MmUHL1pUWmdywIxfTxztU4RfbvFDfmNWDkfhlDNKkluVXaV57+gog+q4zH99KsjDXPsQJtaw
0uRNs/nXdsGqT+WaKJJeDfnLllOKVlAT4S32Lfy+io7FEHEbTbWTKccIvTzA8IpxzmXR6epotZmA
LfGVBqrazVUEItTsoIZNbfTCH9hLdyjqQk3TJ7WB1VdqXedhy1u8DhSR8QyU5mb0UDwI6+iMR65p
Q0+PKSuvdIb6wV4+G0kx8MJfShE2hMMCXxyI66YKaJ2CcCFAA4igL3Q9RRMS2GeEQGyDDGYZhyji
O2AUbWMBntIOSzpbRJJ+GKAh2nYpi2svzHpKVmXW4VLxcX42JgSb9Lvs54n1xFmjOoBnzn133VnY
PlwP7ZxusiyZAd2cU3RahA2h/jpScKGk0ye7951R8F+fonPLxfP933G6Mfnlr8OWTgSEiq9dJ33D
4v/+Q3XfwSR7dOlMj/zVkw8luWVHm0ueb2ORqqNjRedldVJLQl6UFV045WCDH9kh5TBWqqt1JkZn
PEMmko3TbOvo5r70gfGrPDjI900yj2f9f00CvbUCBfnfKX13NFLMwklYObD5J0NmI9UG1tTn+c+j
+R24beuBsXnkTKprMBSwN1z3MIX1bVv/3zNAIOqEMA3Z/ZdoOrk55Sw6M+0siql96WaZRXJpXFWF
luL0kPuQ00noojjDicubjQFeRFk30EkY5MkqhKGMwrg+8HTo6xnCh65npdNpd83++MJK+Xoc3deB
IPOJ/CVhl15U9DZVvBprNsdrwEr7uBdSsSvsyi8kgQomE2adZwQNfWo78eO1lyU5Y3BS5pSEECEs
E3Y/VYJsNFp5kzMoAh/SR/XdvhsdgAHmO66hHgGIKsOitIyDQR1JaBjhdyMRmYK6XHbiznVDw6bx
IjUdIzn+ckZUyiFkUCqK2rCgGBJ86ItzhNkMPMJ9gChQcqK3nZg5FHVfC9ad+J3iKWwEUtNQSdkF
oRiSFWuFMayu5ChDEi0DaPbtlFKNp2O9zM94fNopL+H2MueoZP+Io+kzglhJ4uqopFbBMzQlBTbQ
sfdD7668s6uFCq3d2TBoTwIqvILqZnAjQ/GkO36jF4tcax7YQI36MeN/IK8toE+Xwe8T4VHUqPaI
wgDMGwWFBj0ySIHhG9rNgldpSMPeMKtkNARn86U22n40zWABzc3azTqkvZyDgbHTI1KaTPH5oSar
ijrQok4zv3KF38eRwzZrqYAOnQnA0Ers2fbDUAJXT2Xwm7vsOPwW8Iu03J19UUnhhzUWsJ8cEq0N
zSUbKqRQSJkajrODU6eSxUbGdSuROBJUaIfWflj3vYi1I61FjyhFkXfVESc+11b8V8MlCduQQBPg
DhXSVwDh13pnzLbGyldYnlnU67C7YhPiJbJ1YVfVDC40/NS1/cSed8LEV1/hmcVq7djCr6gXQTk5
e9d3gONf2tVkCA9X5qu4bMoxLLH2wzjqaPOQ9fr4yo32TefzuctS7On0LIVJcGXWVFQBxLDyW25U
7qnDQyeTCe6e3ygWlsf0t04Cdu2JjERUnvqp+aGAgKMSYU6nUYDZG8ai15H2JY9q7mkMNqLWbUHw
tJtH+wF5KWm2mj2r3M/TU9KbAC+vzuwjU2VxDiBHSQ3fHU0pXmH3ne4mrBuWWg3yaaJShtOaIX7S
naGAqmuueXEm/JSIEWq+8LcjrlaXMDaiP1+qeYPdMyijI8SzW0QKi8X25vZDxA0o5by3nv1IF29O
Ifle4rFQyx3QPSCzfszJ2R2D+0gqEM+yXN96zuO8IgqRDQYBrxCNe1zKu+7IYiF3z+nQf5x8NrTR
kVF6NdxFcwjhso+vYAkIpwX9PKrYvRQf+/ORSzIQlPqAv9KqzZeti8RdskOVT9T1mgWe+f6JrSvl
T/XqwuW3MQJCA4XxkZ+kIuDso+1Oa4jAHFZ/O/FSK1eMzQiV5WJ0No8hq45/oV/CSNiUC8Fj+eKZ
kmUTDqJO8lGeRV/Z0A0ARQSsUCsURr5xiJHxILgoCfI2wEykxVVgEt6KR2PV4e9GaLQ/kA+svZsJ
+/mDWNcesxiXQNngZ6LfHgbRqeSoWe/OpuzDedqXuGpQbztZ/MPz7K3W7zIimxoM193h1B3cWDDT
WT629NC9XGWAjSpqrS3LGNmTomNLgzADJ+0m26H2+9CoRFXgWC9udTyLJPLCKzvvqL4h9M0T3EbM
GimrM+KXXYweLHXbcEH++RnlMc0wQRkzAMS3tm5dn6RscN2uIqOn6vs8dXCw4WCcCIxqgU/LTr4S
1NOhs1KwYMQiQ3JA8kwJ4mAb/sX0RIqpub1I/k5PaM44IUOf8ldqos/4AQRkt+fBwWnlqyqydxGX
ya/utwQwr0lsv4LfPP/e3GLM8L/WTa2Ra3v6STf9wzN+fM0/amIeTPhkXFvmOaIztjLXm+rQ8a9e
aKc2TTMPQY+SI+925LREObxYFYMjsMoBXE+hJdzjnFC1K+gAIA2eWiTqATwSvCoHSHHe++GbXNKi
AXqJMEwksK8nWNbEVGYzGm4u71JtgXGwvMlSTJTJp6ozZZ1s4+721jv3KvQ+c8Q5Z0prQmPCpnrJ
Dt7CUK6HbhHNT7nbkZE3p+uu9XeacYZTB6TmloCzTi2MgS7YwzMwBhrEGMkoPk1wnbQTKAfE3fGS
ajPbFThak9hIBgm6H0iFuFyJBtsELk4eGhxsYSifRFdYBfgZmw8Pmr4cU4aVyQy33fwtd6bfh5mn
C2BnZ7g4l4/HWrwO92U2X4RGUc49wLlVYSrzi4wOj+JttCa+7OhE3dyUshT1MW/dmyQYs/AjcMIH
863N26W50jvcMy/32UIReNGpToNJxzMsOqwKh0WSVsDhaJwtLGIhyv54ebMua+gr+MjK0xu00/LC
ujfaKWDGZqjaQ1y42+KYpkyk85VwvsYLgy2hwliuXm9lfO2GHmpmfO1d9vCqsiRleF8u1Kr1lvYp
qWKQ/5UlJqrkWarhUSuY8cK/37FlFCAyxlE9jLpQXj01/2pZe27JtRfN1oAinrXc6y1wkJOTJ5zV
X4SHPwYQ+Aefu51c1RaDC4ri5dYY67zNYWnzKMKpOmQrVS3c5zuDJgk5Unui0sd4w1fAHmIkDm+O
Xpdirph+O0bPdFiBJdQL8VZJqOHxZ937FTxvp2ZKGzBF4aeYYAG5sN2Ba7dSMTvi+md7FGw1510j
Iv6283DSMRc7V7r559EfZKlZfiUMZ865HbXn/C0ipIsHWSbkSXhl68Z1AcdI6DMBaBk+Irr6JEek
zVkCUswZLuSu1qVkbVL1s+5QaYk6pIrxZ+/4dg4osEblBkzQ7HQnWjbrpGYUI6ufu0eqkyeTB0mF
jF6SZBSn14oWN3+CYibzpWo0Wy3JP1YqX2WdAhQQ2qFQ5ru0VmIzDShxA1UBGrFtgcmo+Vg5FfiB
TR4dGWnfw9ugx9E+lEBJHKKbOTIXaCcf4Z50831cZfM4ubzUXekqj45BcA6zAH0Vqd9MmKesqMUg
Ll87jyTMLsf08WBCd1t/aeuhyjTbKnCX/Ff/AsnzqmcdS68D8fAcxPjSKkeIhbO9nOT6SLQ1unZI
yoBjMxSBrBJ1GJs9cAiTHxYE7NbooLI18f2W4dX4mISDbjjsQjCWIiEnykQJM1fRRwh/PTd8S1qy
g2PCjVrFRkgyhPnhTKHa5Wbx/UzNg0lTcmuSxo4RRxJKzVfm9xAXZXLPvUJO1ElwxQ6toGAG7wW4
WyVMyOelZrZPuFOifHNMdHC7kHB7LB/b5tNFwus5Jk2dX5gWXDg+/AjRIEaeM2EGtPJMjNNF4Oou
bi2ebxly2JNU0wB8xsaV9Iq4iN4riJVk5dQrwffrFwmh257r2fZSoRtidROdbq44n4Vg4GTNq+DG
VCwJaydY1jZywNDLqjeEMxbAex/geoflsqLJHILOOq7PZAp7Km7L7484FViilyTJjTk6qB8Me/Oa
aag//ex4oBKpWLNZV61efDZik3LA2W1wtTwOIU2ulcpunWReCpyk6xpXItmT1kPT/BadBVH+QTIh
GvSEh6vFw1D8jbVFGCzU9nSsBB8sHZReqfa85X02kpcQMYPeSNWuTd7+IlcX04SX2zyB3rI1fIJ0
2sNbdt1ANfyZGBQQHg9wd7OCOp03IfzQ3t28vR4GIQtmJ4VoSq42nqW4u+w1ZaS02DL6NzitgDCl
AcBJ1Ckn9xdZdPJGvys6yuEEk5YuVRP4l368EtWEKJI0SvjJxEuP8rYup0NL5KLdozvbef1u3bvl
nRMj7A3UNSYi6gkrBQJ7phrnq8SbwmRMYdRgS/vZZ330wic35moI5qKjSwJ+Rk9/de7S4zM7I/Hi
jaepZq0c8RFGQq/alDJuFymxIEwI1xR7EatqC6kXxwWvWdaGuIE2vjtDAtOkajxKvQ1gngzAevBi
J30jy2MMFBeyYTSBEji7sJZX7yNeqwJ1MPlc9cPcnnM8qHCbKOtyEzpX0qlNOktDINkqA67ey89J
OuPtqCDPCEz0JtGT1e/Y4Vf9D9wQMUXgraK3abVMrn4DEYaPZOW15nh7ZX6x7IIJJ9mouvRvQGSK
g9/GGZriUAs4GCziIUuhEMBUHjemwfXxL8pCVcdZu744ZJahoAkOtBA/UtcFHGPuDPKkpmtUxjin
TZtsLHSPldgs94HScsHrmAK3u7/HzkxqbkYjqgNrf6r+wUK67zv/kYu4eMOrbAg+IHZMV5rdnShf
OCJGCfFiI3EYDJJIZTrYhVY6/B9tFmoCG1/KKgzm5C1ms/cnFELrMcaWLD/w/XrOZXC7OXHPu8gA
K84SfwFIlf9OW7bL4Yo9Q2UuJ5shduH/DH/yb85PHY48Bn8ewvJvNv1TDNVyJoTGwDpmaDHoEJE/
AeG2/hU5cg1NFmtIPjKrtRtfOaFMc+QERW0wh9r0z/dWqX+e9ijeXt1pAgyNC9XKnrzJHTW/Ox19
y5CB2MXbsyZePjySUfVbAgkzXMLOJQUmJTvYrZ8iWO7r+hGXH2zgz5+UVDzsc/TZ+wNOPU1x9NmV
3FJnaFwZzvzivYIkaxN61EAKx/Gf8S1lw01/l+VziSDM/pSe2e5d60XqDQtma+RB8Kl+hQoLEleN
hpklySOO5N7N0hzPsW+UNPnTRiDHR5qGj32azeMUWeQ8swBCwsPJjI6aZARedeqe2FI7+q9Lb2LN
4Pogde7T3xZQn7U/2sovExHfcRdLf5VFzvV+pMh7vJ6xJn1gTLD3x95nWodrm/ezkMhMRA7TxF5B
rm7sMWTHNVV4grZh50IxrpJ6Tw7867Fi4pyRqsGv8p2Tg0m8+HpdCRYA50X5eyoLaJOLoJOvMdjD
QrUF7Ao0zNf3DdNNDEXJBgi5InumPK0yHC8ZVHmoYmqzkECaeLENfgEGv8zvlO3KZOgZ1oUhZB0V
hioanPToB0x3LEDLigBRz3QWSlLUPxc5V299es3nsqUGeVhQqIGeI2MUZLzNxlfw2Cdt3nAdoqry
NgoAN8260peThG2G+suXXrDuxZyZxXsAPPHZUVbhzKiHptEc2SMzzIXErL+AYaPDwgK9Wo7ebY4V
p21sCpoRTCwkBOo+ILv//TDs44g0sDyYRlIrFLGEbAkVjFIwJ9y+5fy6TTT84UyPXU4dVmbhWzhi
rh4P3zGtlA2VO/EvdZAiVvA+IZhFHpOxdxR8uVzghghfEax23IentLhhhEVEgvmR9eXCv6NJhVYY
MJG5kuL6wyYGZpxjvT1eUiEuIs7BjR01uMsNGqBaK8gLcALZc+IT6pYZtZdvBhp7FtfvDjnps9/b
Zzt7qHFgPo7LH5rWCeHyXwiEtmLSmpcoTaA2/TGNGyx10NcPT0ZzxjbcKertYAQ/8a1/r62HwBBT
c0/8F2T0fqb2n+KeB1+VEU+g61o1CGUY8ya0J+zYaQzqr8ekT1wVAOQ9IKOpbc3LW04QD84mqzy+
fMiEiU80RqIwn1V1CKtr7pZtsCfFg8Gg6gFSNkEAKdkur2Vw8+BSf4jcn/zlorxP8A+Wd2J8cZaA
f1Slb3q2QbIozjR+sS0oVbAPPgDBJ4y7mklXdrdEvcinNuInoJNrwj2vrb+rx+yPPnhk7VXYuDH4
q1tGqMAo4lXETwaCK9sqAp6/NI9/0tgyU4eRbzjyA1mkv0ghGvh4lhEiX6yy/qKawCmjSQNDReea
cRZTySGVkD4p5WqyeJJq1hn8FoXRzqw+zQM2hLuw3ahJBVY5hshocVhEKOMbW44cQhFFLFbcEVRz
JHOxHw+sz7y8gzKdXlP3p7wlinANmI+8gJrxQhq2XmT0bfOncm1x3ddg622bh8IZvbzt9AyN8cJx
Gj1fzPSNSRHX/+fKSP50eDOjsXGzps/VjHYqGWNsNdrq4jZtFH4XY3Mhc/PaVOIzl205eF7S6aDl
XrFwRpLxNDCho8JXDQA3qaMs72V6Ml1lx5Yv8Z4HBALfEZ4ULeVuXG09XPQcm9/Gto/2HAorpfsm
74KZgAjh3lwPM29el5gi9X+/lGYrFOPLE8vmyCCEg34rBfqzWnaHPIpBKmQN3Kau3RqVi4ry+Tvb
NuzVc4WxAVeU9RUNu8JzfkRXe6xlCN1QcJUJvbo6/8HBzVcoQtQu804noy+w9uFaWOVIffxBeKUk
AAuX0t3tgxuAzI44iY5LkiShhD9qAEWZfbFk2lxLJKShrh+OmGGN168OfqOHSM1YBr3n+27g6fQD
+r6rRLJfj5sOIaK8Ln6xU8WPvO86mh+JhEAdDsxPgO7GUP0pubxFgb58Z6DL6JhGWUx61rOknLUV
R6FfY7bFhViDN353785nBZVuhUdHpJapNmsMbyRNykDGWpHa4NKsfIZw8wtPpXFExb2vOAkMk0tw
RQ48NeDprU1LjUWVi532pTYamHDsurRdbOyemGgkM/kX7AmZB/RM2vnptlBx7OVpqiBixRgqI4gu
mMCJ7Ksk3vIpIbZDDoTFFTcPJyY38PAh9gq8tbfD53OdkYJieLZx+6xNpI89xw/FWkpnaVBncagt
1Wba8UwAGMB4FaL+IGYDVRwMx6fumRCI1KYr+9l6nyOeaKpOYXEcTa3nNyK67zKV+77wstbMxsKW
cLXEtYIg1frWesWqPzXjQhHPR4YAF2jS4OMD871Ry+zRhVausSpbXgeX/Iu2dJZlQYR3rb10i9zb
X+DSALXrmt2gDix6wC1c5+MnD2Bi/oF0R8xCQ13F2hlpyxkvZ6jedLEk7yXmsgTL842+bwQvXdoo
CBYSkBjdZCQQYlgTNAEcKEcqYczX8IA0IS5nVqeeYTUB+Vh47hD2ycOuLKe6cDXwUCS5qdF0l+WU
mSlerWpWZKlor67tfYSdw96ltZq+MfO+dmjdRgElcpA1+BPrvqxYixBLnkcIh0bRlAWgQvobXCgE
WefZ+em25Sa2ehHM7QwFKjw46nEkTlg4jkf0HU0W2YWGh38S1DHoa4rERU7869BSS0RXdV76qzCM
hO1TGHUgtgGpsXOWzifSGRDdoR8bJsXbSZ6hPQeHpf5gVb3QAmKggdopOdTHyx1rrBOJ6j8bNp5i
2yr+kte1kX40B2w8LOQwAG8HUS7c4rO/uFAcqUlUdq8IRA8GLXWLp6CIy4C7UMmcRdmNYcTb3c3n
1oaB0d2+6CbVoItbNtjtudQ5RtlFCxMHLfOzyNYXFuiMr0ZtrIk9sSb5qBYCGFbmTDGEud27peis
qO/QMrSA5D45T/UVnVGhZy8iCT3o87aWJ+zHadvEguOKqsgBWnOVovkMVMzRCfYvdolvyjXH/qK1
KMSUCqQlU8kPwDiWjC0CsWlszPhVznJW3Vh9ifoPx5ooxPpZ3iGun1cqV04hQl5qponCyhyQtdh+
hBvV4zHc/BxiRP1ojAuz1bN/uCIoykWIqJ9d7JcBuPCeQiWqF7ucagdudZyIdArB/z5Q0vni5W/w
SI5eKsWJdW/LNoiKmPbiluvC4T1vIRdctxIbaKhoLXGXXs4fDedRtgqiO0QOHuBI+hU1B1vQle/j
b/pEOpOz501s2wjJbsit2Yt/nmD08nuW4FTRjRpaW8Tg0tv0sUbB5wUuLzlZIufS2/F5axphYmoz
Hl5ECU6ppv9RWYcZ7TbOKd3bC5E6J3O6qxEKehpPpBpppuc5QAb0QdQHAS/xoZK5YGdBC8HZWLGt
+7FhAxgPboAGLqRwkkeK/7B/gGz3roc8PcuPXDQLjKInOnT0+Pq9HiwcNzk6tqK+9UYhOsSgK+LB
Bd01/bViVCBXYDRwsixLYmwPCPZ6GZLYlOX4uavfBSIfQHuF9VSWVatqtm+yHLLxHqk/6rn2Mf8g
AkBEdFKttM2GNmENQPi1qwZYKK6pQtzh5eHaskiw2m55nJkHg6DnpZEhK/lOJa7wdQxWYVpfTJMR
RBl/YuAFnyYwZj5jmdFjEWmu+lNB2vPAw+BCYK09gDMQmbIDAqzoxSwuQiQjNS/47LK+Nx8+u1S/
e5Dtk3uh61DOMjA2bh+pYVeep2l4MjDK7EczxGHND3qkKJGb6bKage/AD91yzvupV5qrnk/bbfCi
xESe/LZuORrKVpY/c4tCXNm2bR3yER0penOsRv1LqyhhrUMnMUQLeVpEoXnumK986IrSy3VAAyn+
LpIeNSgr5HYHjjpefS79SEIMWNTxwujReQ7Hs2QvNwQ5sUIQ/8HHhqK6J7kgtglsAqO7wPrdxAng
35zTge/cwdd3Zx9kQGZnu+q5A8PBPJIUcYElq5v4/c1xZfa4fvVJB5aFBZDfj4YSRS9+X0YLQsYK
Pe9n4nI8Vt8wKBq56numHJuk1A7DMkP79ozI95dGyOqdNjPI9+AAM4CVgZSahP76GxRC2j+ciogP
znMSyCHeiPzonebfNKHGplpYNgU7qa1g0pJ0hkGFQMAgo0AZRRqZsa0NASbKu/Gc04PgtRVfW4xD
UYX3ATjfj/60N4YyW+3PlKGBcpxAVtKqWButcK7BU2aFU7LoBu6EAoOE+RWRtHoj3upnTCeoajg3
TSpp6/EU1x9I2IRJB65SEJMSpYByxy45HzeWl0McOo3CUBnEjFDkQgmNTE3e1HXzfEafb9n9sOt8
Sdvd+23IpwaEfh50S4JvZNFO4hTH5+IMCH13Yu+S1MMbMe4iCy3BEJZ/mRxOIatOWbgOl+uvMCE6
09rmoEEMtUzlH2UjJovx1Q5XV7IidU7gF1p4ceDXpHUB3oKkB+Z1V9Q6MtgBFOxYrXC1UY+TP5HO
8ALqG5VsR4prQhsIgBTcx70DN3Lu0R6uZ1hax4MVT+fPYdiq86usQkFPMmmWCcv85vHARK7jmMB3
TDfABdw1CbZt1D4jkDaqKXjvzJTHXzeE4kRA/F3lHo3FvoKvpZsQ0g4dRpzEePsR/VA4A0+ZWUx4
vs68+EonCXq9CX4EccfRMm+KuGGm1bUSGBJLcTXMY7ivAk8OiNmT164jUerrWG05j0EsCp7JWGUu
hueh5bOqYuU5Z1MVSgc4ksxYF6JszENfBWBn7IrHXfmjM+csRB1cBmzuY6fBdz/iLhMyq/uy7P+k
JYQDoSLt/+TGUr2wRCLdaN/8t0CAJNtwkd8XG6TgznCMf91JyqS0mn6GpIY4IilgqN9h/ugB+YmN
x+Scgzuf2WxJemWqPn43T+/EmcJ6PLp8lp5MFAch55Z9MQJUstHz1kZlaNDg9HbQIah/7EwzzCpK
GFZhtbiL/kQfQAISyiejM2sdFybaNmkBiplO+pD8DfTpRrjKvXnsQVzwaAZ7YA60zC8Pc4LPqJ9f
Gaow3nL9kxcq7qwtmLx5sW1OVKCmaQs/8YT1cSW+iMQiAaTdDZ3KAiUvfhQw/T+bztmccMfz9e6I
4nFsDDuyAEgTgbgocj3X4/hIR2a8EcxmnVKPGS0F21EpS3STVHhr2DGoSFSFQssCqzSMsTxSpmSR
9yY0o/NjLY/O1PphuLselj603vOsSSCnAmCKkrdPt6jC0oouTFXzOgHTDZVOc8fCZtcwgNVl0lrH
sPrskA/tm2S4BPPNBnKPCvVsaGibIyJBdS4OuvAqFrET7UnkxKLbNE7NTiCjRrNS9fCKx1mgHttk
bYLjrC9h7g6hsXi37I+sJ8N1zhiGGKJXbNm6//RVi1tFJDcRro3L1VtkA/wdF+3QA7JnuoP4oeXO
kR0VxTs26gWE+PpPWanHxMM7RuhmhzxlD4LWvRTuxW3tHoqi9sXVQVVIrAwfPS8TOzoU67YnRxpK
tB+e6fkE8+/VRmvxbhf6KLn7h+PB55aVTsDIpIhxOgkIA9Aedli0UUwfxCjt8BwR5JdSAyYe5MB0
MWzh0IbIlTgg3OkpMnAlMTd4gF56jTj+B8SdetYT19i+eNDyLYKniQLgTcYhQImZBKUlPOpwbsQY
2aoB8wr2Txlpvb7DyZfa8GNmizwh6XZAZZjbZNtPZKjJGXo+fFPmbA9a6IoQwAj7a+NSvX6vK5As
j3O5o6MEvZkhMR/ggHvgbD09DkCOz/PjP8dYcymYUppV0cDc4yElhbGWZwEu9EDt5E0YLB0M1EaQ
bxyLT85QA1VOJeOX8o1yTf7OPKoLSgXHe8C4s0/Hu8vwqOEcZKVRJLutBJTRkjUOuVvaMzDM/JiQ
q2kGfyT5VhiyOBxWwZNdtxVE7xSGZUGrUPnkUhiT0LPVYgW9updVjqj0qWeD3do9KPayKRdYNNzr
zxSibLmEtL4ZfQmH5ZqmRC2R9ADftjWgRPiNr5s6vex/KpQ8xJ8oiqbYkBMpEEIgS8G3/0kzWoNx
7qdCcJwTxYN8glvLq7/iqCN8Q/7Mb6mbF+sPHPNDyMw2aqJSKlmGyGXOcXv2ter8aZ7XrQ0a9JUK
4IzbML4r3osxUK/KZIePPKVKK6a269t15El7y0rAa8Vwbjpjgl4DNjWWr5lzno7ReGFaWxvqjpke
V/lJTiGMwQysZVdUQ5mmOZMwaFCveQ5b3FlVls3PV5nRf7oSLmbNNZ+5Ax4LWdmjNDILXgWHI3h/
btwLJ42Na3ZLnZmoe/XtX83lrIOinqmc3Jl+MAtxlGfjuQitxBXeKG0pRFcv/Wnqe09XLx/w/WvF
sFES6+i9SvO3CIUBQuMF4NFVq18/Ew6eDFqxAmEZaHVGfOoPvUrFgprBNjDeb2s02/W6atBH3y7U
Qam/x4JjyWhd/c1FI5gN2J1rgaMc+l40cpyA9DpEXgu9M4OQnAfLHkCPS9nYVh8ahTt2WuQwDl0J
WOGyAHPkE0Xtc7iOE87nw4G0N8yx3MOW/jtHU96zB/VGALaZ71GR8iggxTMu1B0Aj/nBrkA6THrV
l/HPEoDM8FttWEjhXg5VviT0XMvN5hJvHVPXx3rFt4QDptDAOKvxao7DcByHZ0av9TMpSeCqCyNA
r1wLeFT/mZ1hS3x5h7YVl49nW4O0MfpoET2wxQKY1yT/IPMmFm4K70pbE/gk+xmhZllmsqJA9bin
wO4uwC/E3fujMZ9Of4gY5vZZpK+hNIQFU9DsKrxxotZAN65gTN35611u34pT6qkHtg/hkle9pMi1
bA9lMlO0DnmS8a/Tn5OAYQOTNB6ZXgYm4kGzcxkyWxkcHBeD4Q072Wey9CwSX6WVkeu1QaPt6Nsr
d+fRyxdgzfsm7adqljKYn4vCr3lq17A9eg850eGjN+EcGQBunVanA8oXUdSDrfGHVbDsIBjwuG3Y
hQYXB8OwVyZ4cy4ZRHEtEgXffXan6JDEujjlhofJj2P89PeV8/G7QTlp/vkpm0GlbIa2O+R+Y/zD
YUYAa2lI0Rc5F/s6BZ30zeRbcwYstpj2QKWEkEMDSQO5g7d5myiAzsEtFiEbxuWib75jn3lB9rcl
Zo/HtdzScXHdDI3VqnaPwfvooPppDtkbG2mppBSI9aUixVWCjbqIWaGgMDBlBkZfK+ECfGpLxGRv
UFAeepQlv3e4CoRKc1hA3V/ZZg2CXNyY8OOksAeQqpkDEb2DUEPDth8gNfodHvYSRjHNPWKv4Wod
E2eF8ao/9oHC3Uy50wMjSdjYfJToOJUSAoge5NcAbxUaTSZ2Lto2g/fkvaU+9siuP53bOHVKJBWz
vOXqSKNmJaBRS9nCoeEXWSyVgceAFskXgCzMEDCYLANVjP8rIzYqlyLBZSRVN6W94QQPgLoizMPu
8Gj/4XD0DhKucMLGyI5Qm9XfOQSUAXAqJPcUz852peMP5TSXIy8n5985ZQWo28bfbGjH2gF1VyDN
dw9v55BXvian9xkL5b8hM00QdAozATIu1rYDR34xH2i9gIiBE8k7IniaBhJs5x3BN05QStXsHxwf
atWsM9npLnGuJIA8kkhxKJHFYnm8Rr9kTMNa9zbkljRif+tIRV378BXFZbHP3PHl50CzywKTYvaM
NDpkkCTGkVdlp3JZIAjNtuhCEuToABjhDs+HK0yu2Cl0iahBo4AHOlX4yBh9MpDv2QcS667trSYE
Ivsm+/EJKyviyKUuboZTSa+L7ZazjyDC2OANx4ZSEsNH1WwQPSVbOjG7V90RF4CCU1DZei5+GP7V
9NpbVIeif4ejl10MjQe+nTr8U9RS0my0enIilzfF9asYnBELjgIH/SljGhIHA+Yu+L+ieLNLoXe7
4VdJOqJmbj7H6XJGI7+jZ4mV2bdHj3sSVZAoJt/OdRpcpmlsgRiHUVxMJK6rJYUWt1v7T+QqedA2
w5/g7Gi8TebcrMcb4NhBdWkobG56+GiU8Tk4JNaQ097jOJm78GNj4NlB8FapNqYQAulCjBboNY8N
4Or9IvyQsYpJAaAQuXIJAWlsOdfuZmRdpyYGRqqXAnqZ1pwAGxwCSlqgoykDJzFea9hywseBFlsf
/Hif+4xhCrKv1VgZ3jIr0JOn7/cjhvCRQrSk+55ikXNs4bWkz+nU6WOJa6bDiUfaa1PlQxnPpLd+
eAcLH0MtDRFwnsM8qW5SBaJUEkfiDzvdyhiPG8HCQ9zVD55gqht3AWPGIAsnakIdqyVjQ5FGeT4o
UA1kaA16AhaLi/oqxkyJiLAGQ/MKGK22XTXZyGNAt4GXU5XBfVp5sOzzWoMHycl/2VKnO32UXhL4
42Iw2XSwonPFHZcRy9DXkOW924lJc4d900sdkF9TXbhjGQOteWSIPLzc3BtiETqPHUDzuiFU9+Rr
uCAu2h9fFIAk7aznnLPeR74tinpVjKiDA7c8KhqH0hITogERlcaFcmlnT8DvVJcQ5+vgcRgBYlt6
xIfWGqRrYkAvXG5dyv2puf8sGEM7/x6Ph1/B6iFdIdvoEzi6CLB7sWo/XQSuRrcLIAequHDTZpHu
X8ebr34JZKX1NtE4Uz0c+BvHZQr95ZWN950elXIeuS+AiLPZVlEz/eNI6GYADZ0jKJLeL4tzGnag
UrM6TFeQ8HTGOYdUh1b0P53UGwO3jJjNMMJiX/URrDTGdzqbVxK5/JCtHeYUd6RlGUC6gNVGzYz5
7bFwei0JfHLn2DV2+SmQ7C+9Q7Gxz3b3+S4zj2U6YR2PKVbEovKoRlzrU991DprBV5zdDIJ9SSlj
JaNxR/sn09wG5zHagvO9XmKjwViPnrnBqXcEqfbXCshh/RPeiakaRlqsPIi5JXrkd01vXQsE8tkM
qNl98Cq5HrEYgUySG07fLfE2gHNNhIEXYhlSb3ydNFpdFqB+NMcLktqfOZX2xSxtZCr/VAPczYmG
9DZV3odUcO+KHxqkC72tB3hcJmr1qvw2Dl6HeiHTAeNee/AqHUzxz2nUHPk7M8FcYLP9EQoPA+4d
hhkVzE8cZXdkM0CT4FMu9BjHH0KVdd57gOrDrf2qMV8gRqbqMYq49N55ge5e0reaLcdKYPwsBMa1
hqHVjYnFW4nZZ2h/NFHi3V/ny3gONqXTwDukmBk2/zDs/6iLeQtKqpIhI7LsrNT7kBF1i32iWwvB
InF7O96sE05nwA/ybY5nGf3aI/p2Cw3Q+D7dVPQwHFir2b0VNaop8NAqDX3hTXFw+QporcEmxXVO
DSq6ba6Youp66CQimMogi+uGNXxNcssMTHnEWJ15ufcJmj9GAFyOIIfiihGiA1w+sQAaKMX9fdYm
yttrO2ayfS7lkJSKBqUkyxzB2WnBNoTQhuYNDY2rhGgsEApjNiPBmKrY8BW+Lddxeh1P1j4X/Mba
FZlJmdcugPz2nUNDr1tOwEkQ+IwSlemYvoJgt5nYAFl/PdYCDBCjumvuCVxOMR18AeUaQew0hDQb
aaLkfJSV28Nz+bB7Vl3VGHoW8ZMAUepQPe17AbPabl8KrAfAhZPpv9Ah7CpjIbbEIFdO1k+MJuHX
4JZehIJ0BWF8VrXhEmh7OXpJ2b8LvUPK26pnPgB/2QfjoK3gtuLlGQTXDpqa0kBeq5jPlObklR47
NbgCWpbnB2AMc7uvo8PF2/w8+gx2/qLbKtPOwcFDgHpQm6b0V6vYIn/XvyVUnMQxRFRqrx8mYEO8
X5Uk/1Rt7VXA9NSGDBB8smyZhhP9fRp5krje8JyZlDVACu3orUjay8RmNf9pkyyk+AWMH3eToTCx
cdTDGIpU+oYvjeLHHorIZFHVvEv1GaXsCN412oPR4c6OfKzDRW0J4cZFeM5qY01Xfb03JwuO2oKe
g658cTpG0YY0cya0WT2VqayD5Oawh71O9SB0p/Dbs5WrOfImMhHv1XRCtg7+ARJ5RgaFy46NlK2J
wnMP601V49ZcqBwUQAB76FzOzLyhluAGK1/svJaigyotj6iuqM2W3Ww/nQ5iymNCVmPR0i3Hji5f
jyxfAhsaoKAD45IhcLRpny0grdL04wThFYH2oFhsX/URuhyOsB4exksb2kRMvZ9oddrmmCdB5f8a
HyneBkCa8fan91wH+f7jrMqPcvn8uR/zmzvMcCriaPi8K8KX0Eb1Rj72rQ3q8S4XGVf1NvaFNpf6
8NQiZ3p+BRhDDI79ttKtcYQLCfTdz7/q53Hkbe4YDGRNf2iC+uPKIeU+k16Br8oWkIgNdxenU+KB
i9o3GsVUvc7icF5Fms29BRIiJ0b9OnJq4dQOH21fq9nM1i1tkMkSdEMGt7lWf2wnBHqUJJnMusMi
mpuEzHc2We9sGfzhR6TgHadwQ4lmUUB82iVirHyp5DYxji3BKl7cYszCTKSAflBMMi5nQZJ1UpN+
lXUvdGqwZ/yNFPGy6Znwa10RHpCN+M2DXBIUMkiq3cUMgQMf9YfIDHnIGl0c4rXn5yW7gQcNTtvy
hUfunRobZIYnR61rCQCGtO0/5JhemN6aswQ4ZzsTlrBD3iX4VO8hiNbtIQNmPKKyQek1jLXYZf6L
WpX41h1GpGNRuw3RnUxMqaL1r1Svx8ikJfT/Hi/fJMGiNiHGc8s7S6LFmQAlJ6foxYR0wj2U0NO5
jGsZK/QVagzdvJxnaDdWiM31jqngHa+MZkx4oAMPCJlZCtepu+3WKGNtoyssCptKZduaWCKvR+GB
0SlNCUvvR5JFuNQoRHqjcBhFLhClQhayYyQwsdguwGMZ4KqKJzt48SiTTjyIEKYNww+1343MIdTf
WxTSqJ8qq5NDXhzOG0O/52QfyN6f4cbzUXzBc1C9mFjeQtoSiip2vPyS8NYTJWyLFR0hO+1b876y
eaV06G+B2aSZSR+qwkzeO5CofNWrkDf4sC6Fj5o5SUKGEXRWNoE1dUZBHDuMc/3dcQvhTuSNRTJW
6gcT/m3IJypoGkXtG2nQ6IUMsdwQHNmvMs/1VXIuAgELc6z6lpa604uZ7VkhZwHNpZdVnxX7w7EJ
DDmiecP+2VKflRv4xwUc7PK706g2FwQTpUVVUrJLYxB9ZQnW2+FFggXhR9MtpdGsoOkG1abGSV8K
OmxUDwzSN3J+HBzJbvT4NA0p6BdKDubauk952tVcwJqLQo2tciEO2nmf/BGjdxT1E88NdxJ9LVCs
+2oZ4r69h2fidRZ9hLbVj3lERPeOCzcV3yV48vcsvUDSE1IXQZ/ZhjaYivcTlXVIYUxyYxr3Di7L
5ue3Z1KYPTnyeoQJeW6rQBle6QZ+QUUN6POlhd9gLutiSNmSeUSMDI3cH/5wd2ByadxEqDRlKMl+
K/8gDZSoGXDfwnO3GY6sMYviqgyZ1K+TELSMh4viSaJEzowIr4/Vldsj02alS8vRVQ8s4tR/bAM7
j9wWnenz0q920H1ft4EYzx4UA4evz881IQvYO2xU5InjSFn2OErbcl02foXBwRBLdmPBfGbtLQC5
V5MT5EXYMrwcVhcIXZvEdbHmxsg9xYriQebLX1qUoFermJ5FFn+OmqLK9V2G8YF8MGDEBoXeNS/9
Y8z0rkmd6XubquyL9qOo8GRgd8jGvBIwM+62f3ufsMytFpRCP5n0EoKqMqruS/SaQjA67XDzhBVr
BxdRxLEmK3xE79ml1TPr3wI9tz4THEEaDLp6qVbtTAGe7imdDP7y7bSnSWy9AZSQ//A5lt8KipR7
/RuzQHDLRWcjh0AiKfiL68nzlV2DCRI2NTVcOgVwbudleaRscJTSpexhlBWgEHC2n/JuNH3FAtGW
S5yFaC7wyrMuwlXdYBlHeUZYEQeVE4KSOXKx0H/qveRFJuiaaVdKsUAGXVArCZduXvwR4sO+tRn1
IBXOWV8F+Aq1Cy/XqreVmkLZGVEduQ9L8yXeBEIc1Z5q4K7xnPwO3MiBXGRg211lahmfVaRc2i9C
xIoLQrp1JF8YEz+3Mf8MsUlfCNL1Ul9Kcn02thXvZQxKqKv57RGp+oQ1B90wjiDQSemmqJJRNULt
es3Vp1xOR6ajWnY0KjxKOZvJJuT1RcaNFDitI7Em/9GN5SIaoAn82bnCORBbNwT3ck9aGNb75UQk
peCl2h/rbFx1F7b3Pdm3uHR2ie7c/IkqD63P2jHuf+QH3LY2QkVsBwDQcSKytFso7s5R1ETqqcQK
5BL+MaihaJvKGldOVxhUfaJj5cXrPv1GB2hzvu+JnUW6E8mEiyYdFHB/yt3fbhIrWIH6pnHnBiD/
Z7YjFDSz82cyVbgXLoXYYdYZrgN0dr4fnboA7vFt3TDCTILh6D4mG9lzlt9VbM/5eJqIqSUOG2Zr
LopBh2B9H5hiN5/DD9GtgiizmuAgWXIQRVXpFcRHo8a+DzNB5UfasD8mJ+wnpIM+gcrma300AO+E
RyaTGwNoQwLgjLi7df7pE9UrRuzYhl08h3oUxpz2QkNJe1p7QtqVQaWQPHc1vJkM7fUSnUnj0Vw8
6A/d0dyJJsOicUZKBpQnYrmc/Wt9tXkfYku8Fssw0VzVa+yZlhORd+MZZUcNDh805iP7vnjBGNmA
KCguSh/AgSczvHCe11YLUkXXxi95OUET9mNAZbVr8sZL0U+14fkx8A5lgt778+bFfFf97VcU3ErX
ptEtg1tK0e9qT2dO4fxKow/d8ymrsHfjgnIpy8X/FZm8hJBF9MFWSj3cuPyarTvPrwWHGKJ1ae0U
bDVhuiPUFvyhFARpaiTOdqst1dCG0udEEXit4sGu0eIvDYPiS4+uy3E7FbreiVjvtkn+SlytVNi+
hJOgDQhrOS3VmhheZZ7WfZ0+JCvrGWfcr8Ju6El+fynaurbHn0K6bQdCMfuydBO0vCLFGVvbD7Xj
KOtl3iODWTc2UahwES+IFzt5AmKRako9lND8siPppMcPpoCXEOj+U6iIP8I7AV1jdzBWZOR0CaBF
ECBsRcNDpq3Xms2oCwiNyKRyGR2H2wIJ8yY/ze3gav/JegNyBXN9U5dYX22mxCi8zPrjYTL4/Rhg
25rM+/mWty9hzGM3cX4NH0S8R+YCNh9jL4Z7gHxETVLzVjF/WFFixzIrpz9I12dj8swhI+6hKZ2z
bQXTLgndAF0Iva8/WDJUpeDR61jhkI/dMigvtczK8SiKe6Mhf1xwYWIYbAGFuvP81JYCDJLj+Oh7
D05x75B+AgoE2NqHs/Qa2QmzD3xDal+5D/PgY6yYtqCsP6ixp2nMqt6v28FmYcFuxO7AgNmH8sDb
+f/cTx0++NcqRRjZw8r0vwmzpAwcV0KDwSv3xx0u2pw9wChra0FtDbM1onmFHRmWVQML3qxOgUle
iHi2k9DZMePx+AcikB2Rx/AN23H+DCmXFLSsIhnCT4ar8epO2soDDhA2W5mZseg0tUppIXEoPRUo
lBXShBFU7kfxhJ6gJbLHh4QRZNHe12dsOs++VzA6qVfgBzQQ5mxoBZpsWvrGsaRNsbFriWsh7+6+
aO9IIvoG6wwq/ou+D0S1j+SOOC1HCtBNIhFC8NdjyLIkd4FCCBLbMKRpRYlB/5B/BM+PgI8EpZHa
kaf4tB/j/pcxzx5CSJtDdaCU0ZJm/y4zBnb4M/vigL5afpTnWvSARiy3/71K82/J9sXea71nLah2
WG16ZRpd05Ejt1lCMPb0cSDuGs2p/tEM/p2iK0BBeXZE81DCMbPdYATTopa1lV0EdHXntWbKBXCh
Gtrf8sKKkJrezdkd3ErWt2Dipr1Y/QjP7OBP3DUsWQ6r1n2sV34AqUKrsV0kiAhAAEIiquGKGvVO
CluFJFop2lcUCTbYSXrpmH6RreOIpV17WC+D3dpsdwX38KvAwZ1slfel3QupQ1au74T1towqK4DD
8tgqy+IpiZqkQ1AdJQn4e51cEy757anu/4KMi0RQFSVaEp7pYNV/GQlOVmjUnS686dhncBO9J2ZB
Snwtj9XHxnbz1RIYGB7FGsVk9ySWHL5j9PHpzA++YqjA4Z8D4hipxJ6FqYmtipbWQ0BseKm3iRnz
kchm7y3F8WT+/wcI00aMAxmB6oKunsI/O8ndlHdvAAu+ML9CqRSP9DnnLTn3xWX0Nib38G5G+Ab8
zkVWYXujtFBAi8efrc+rPmJcxVhTvD55sFYI1azJAOLHGDWcbnx7pf1IY6DInTQ1R3qj44FiSEZH
jYMivz/8uc6tNwBCPbQ/ceTvTh+wU+2Pa9KKSK4PRs9jxjYyFRKi+ADUgg6rs4z89VX3fHJWwMLP
9tl8h/Yh88MYXd3YjH08x0UJ2RMYZOb+xpeaKpF1Br3Ayo/xeiCBEEAWl8YWzyp6Tmaek4TctrqM
kDEOig5VLjwhu+1AHg9lH4EorBbyWlZwaAVGd5EBh4Rs0FDrQp+rH62uHD+VUdlcmLI5BNt3l8W+
wh0KXS5/JmQwmGP7LFPcaxYC1LfOBSlDW44LW0I05tUlE9sZ47R0IVEOSmOCqx2iDpBRp1JyUsbC
LPqCS++JOquxxQ1+BWhY2CptDt2RIdOFVyUA2dJetN8sgUK2IcZvIPSXD1rkt576VUxZgo2Yysta
DDjj9f0L04nhfctYShLu3m2XwqlGouxQFgoKxSYHqJiJe45708eNzhh3v2BLjo3DM7WiosOOr4aI
GHKRjC0fgC5qwei6wsIdzySZSigB1DLNR+iwhhrqNRVzEH9TvlrraqgUP72T/3F/3fR7Wp6Ash3i
pPlmPO7P1DEZGSGBhuUBmrXMNrhgihTcVx8nV7ecEwTLqzTxqZlYOGnI6k3RkDU/ht9oTnRWGZmW
6XQHoctPVpiMSmHJLHdlMyr5Z8FINcV1V9k//XLbu45OOPvDdE2mIjg72zlqjyZbNykSXgXkRxhh
Uo5Q2g+DYMnE+AWIDypxuSP5tgguiG8ne6NPM4bByCKh3cTSz5klm4KCdp4kw+gyMgyEL6E16PCZ
8kk8SCb0T16LlGuwrylRguegUsxwYuwa1PGa3EpnP3WC/Jv6c+DLIj+VVzQLQNIgOyeP/MZASs2s
aeNuGkdvhSCmoGBvq+q1OCpgXqF8kzrFQihN1EgXUW2/6KPaPDdO1E18Xwg1Thk2AbocAv81mCBq
gRpIXiIVTIHdhWuPY6nD7Xa4HEOBuL1H23yrf/+WcjIEZDNS5V64SbF/bPrdWA6GzwvmynYnxEiD
BaPwUuVwA+gv+QuBdRYJKRudMg0/PF9nUo6mM/g43xPOjzIlLBei3forTMDrhJyl9BSlO/mYlART
AEwckaAXmNf+CAYLnfr1FccpAnDh/BWsXeQbBgwBxnfmZ2KbssHeDPa2xiYi4OhEOUWu4U2LEBtS
OW3ikzRLQWqGBUrk60q1QzdfwaS6/U1Tn7bk+47fK/csWb60nCqOct0RO28QMtBcz+CvdB4wE0PJ
RqjfPsz7PRA+5xRBF2H2e4IILjXIagwsJiGu3iKTnwyN0InxD0Kx4uHGBDy+meeKYsNbGYxMNydI
WD7nOSL1kEnDok1UnGl0DBKq6pLx3DL98avBBUTEZV49XcTdpLunv+IAY88NglZ0tqvTwOPnxjdr
PnoIy0i1DXnQXyw96LfH4g6iOZm4sTvlNYQ55DKNSTODCE9LIIKPgX4sd/RAGFfIvTDY0ibjc+Yp
HWqZ4t6FbjgZ88EpreavKx75gO1MfsQC6cNf4gsqsN2RdASTVvbsD90JCrQMZiA9TXAbUKWIfck0
TUCtlWyK9mAmHtimFBF/ILNHU4V1PNvNAAwnjAPtSaUZRSuViQY2/+x+ZvGuX/tloUVPOSjQZk4n
q0MlkwXhrJtkxJbdX2YqUXF/RykvwlTZ4KpTJZMOCvZIVcPUVA3i04j3Zvn8clcdUDh4MQDGhe65
CAL8WCTFLG7g0VZ0yi57Y2EOXf5RZqoKk6sA3203Nukk7/psXiDGrVar8puVqs/OB9sFqNufMsLD
7rWTRwHH7ObRQtCk0ZYOCZ5h/3y15qZiAyw/9OS0/iYKK6GC+fUxWzs1WhOmbpK0Hh0RCVPK1WQP
1gmxpAF/5BK5ZuYYd0W8R2+cRgxpb/ODNBQc0cV/3g+LUNb1czZ4gCOZsaocVdNi6nLvz3gtS0iK
NcJ+EDS97uoiHb6gB2fEWst9BvpS4Wbe6fcxEFOjZqhLow1Z9TT5zM4On2UQo+bjenZVpdn7pa20
fn3VOwyzLb0MRc6HgBBOYx5sWLP56+lSUM0HWXo4IFnq+QCEpD3Ucw2lFsBKl3PmAEQUBd9ZaOGD
LSwS4R7dMHUDihfVwEzeY5NSgnATOAZ0qY7WhuOlMB2KOrnF/dji+z1w6iglf9JksgEcMwFOe+rG
wdCP45SN8dRTV5apIqxEqF5vEZdzrV4ufJ0zE1dYaxUGYFRT2eR71lXOkRzr/HMVvC+fr/Sa3OLQ
oecvmLPHeiPtrQY9xBLQjLRp/TNpBHXg3OuI7Jr0qHNptRBj1ju3SjrK6vqe18tDuBmE4Ykl9ePv
mVjflifzdbGSjkhyXFc1x3bMqacgZ9BSxp5Gr8U7uaKQlHvZEOZlPIeNtK+VUA8ugZTNh8Vnbar2
ndnOsZmxbE04/Hn9xV8i9eZIW+4sf5x7YwuaGMJLAnkpxOTCRmdYIzVoWA1dvvR8dxXGWnVTfY8z
7IEVdyFuJhaKCESx4HWRT9dcM9RnOeFaMrs3ylbu0lC8Okh3CqkksbWXyCfKAvVHSzKWsmTZuQGf
bskz8Inl0O0BoUTKJruIqrbVFrMzxEG0/qRqcWDBaE14I0R0UlvVh8EYTfsHv+iFbU2g1leAQCMU
QfqzFAQIDBOxrOGF91rkk1qyKrQF2wB7K3uYngs0MAm6/WrM11+3sZKEQ6qosNYM7R6av1wRA6fQ
WMpvaVXTSn1p3+vFQCuMj4RaCjhSfF2PZlbtWbcSL2KeAgiASu8SNL673C9oN385ezkAHOpqo/h1
HCSSqB3dedoDoVcroI6OJ/ni+nA3Frv5D60QAMxKOnTJwD80KnStU5YvlF1HV+sUH5vbGgyenCeo
mtsEZtuR5SPW5kOnwtPZDcLxuP4+6qpSwkWAatblL9GCarwRdui/227uk6keo6A3BHodZ+DBw1WS
0fkReo2DuCWRlwftGr7o8lsjJNLJrgw9BidRjazUNpuJLm7LKqdSIHDIuQMmSrgnWvxiP+JmC1v8
oTiz644zydePN51TosRYLxtcRuq/rVycLG2unZN2CSQqyDTHdctFQhfwhcW0bbV8XmVWtPz+C05i
GuJyK3tPLvY3WKnoHslxByrFEbRPvmbR/wl14ZqU5x+11xX7s69j0+4cufdltvnLI9Ovw+tCBkji
ZAviOziS+JoSiIXU9GSHytoWclg4HKkHTHSbSoP5am43c9cWOk5QXcMcZu3F+p7xdvbK6KKNF5QR
L4iMgXPiYY2lb4GOCoyjzaj1tKstZ7ccTKsOo2gpfK+7Ig4+BHs7Y6JkZp850NCsccQzmyLECsND
iOL6b+4hLTnHesZoBsYTDItaSvlDJdR6tB+vBXEDArWtRMzXop53cTsF4KwXUaugaCcwrf1KQ5FS
Au90GezghFMrVVvpAbz8zmBqbJXgWPNkt7t3y7WpJzFmpyVBEM6l65QgPCLiaZvrDThHDvOwsPST
WFBovHpisJg3Gv26ldtcZwhpJW3ZUD7jUQeJ1ypzVIqGQd0MDICp3q/hN1sN3MCUFPa1dfSo8H5D
HSwnxflkgGIxGIcgBeLz7TydF9NpUzSCwwfT/HJiBrAzgJZpW1lpV09EY/qIHutS/JcGembFEXYt
9y93Z9L+yKX9JEp+O75rXlpNvOKQOVL4XtyDHrsfD8g83yX+3VQOpiTdg8QsKbrEwSzKqGYjDE35
mCL4ugBA7mAMp38qDSzkXs/eSF0d/lo4GTXQ5a1KTu81pk6ISTnnNx0DC/29yOkQETMjppOqe4eO
cMfq16xOykeRs81ZqpW/Jipdb9lctQ2vFlfDAmKAMF9xc2X3eECgRIJZ7HcFYe/bRrWmdq5IVGWh
7F2nV2kLrMQ3O74nJQRnJim/rGX3tJ46jszeI00th/sP17Qz0kRbYefTuI322pCXNv97eb3nulWf
kFTAmIdv4bd2FYAMvkFt9TVG7kTpRaJAgEmuq2xixxCXE3MEjAeWyc2z9SNHXHtCfhmfHL6LTjnI
k0+GvWPuVLw6J1chuyuo4TUwN490GZrdbpNjbV3hl+iiQxZYaiy3z3r5RNgeJa3JUuBAwilxC3Q/
6nOq6ysMekNutTrZLFuWMdhPCFWLbZwMTb2GVpdkzbuZAiCm3wsmpMRB5FExMwVRP8X8t15EciZc
oHapbS395s8DjTyLuYQ6iWnwE5jn1/D7HBendD8rD33uWOlXkbTEL5DQPMWN1jRyRy7SGIiRIoKB
ThkjRKZj7DH0crSj949cRHfsDfzIPwxhyUfi2rqSci2tW74rmD/XrM/XFkdMvn7y1sr1MHV0pNXI
GKHpTuhNiSygpFGeGH+OldO/Qok69QxrIXpX93SZ7GbdlZ1GsJsbfYNxB+g38uTrw70josnmMysZ
oYjJWxW8rv2txcin+gpkD+K2EE453xndXUhZEILcH67/kXwRNG4Cr1EaAFHVHPmD6UByiCqEwUqW
MLfli9sXQlHTRh2ky1UYbnTr11F3r152lU84dw+lerwoYupuDiiLnMkwF/6wI7U76w3Hy7LXRRVo
P/0c/3Tev6T6XHT1ZPzgWjKrBYijvzmEWV9ImTMwy2OPqcV7zMKboSWJp/eE7Uh1KI7TQBXdZfo1
cc8+Klk4++2zlS2FjE6AT+xFtFEqOf8MVZ8pl3Rbw9MOlvis7Cd6UF7TiaZaoEkPLH4PsavSMnQc
cm7C63hxtfTKWl0DPE7nLVyVfNvAaBYD6zjqdFVFjt50YDuSuxdZurDscrmkinXmIH62yo/GAeVQ
Cq1Jd7iCiFbqS8wgrnDR8urAw+u2DVi9oGYu5ObJ1K9MPLOh+QsGLH9yiSthKM2hUz8EBVXF+Jp0
t7JOQLkNNMbcfUhF50GWFZPxi86qny0koKOldf/lr/YV6QaSizSNveiQlXBrxCM0oq6A62qK84tR
P6omqHk+0Rrf1dGyjQ3YwiUuYA+XLEQSia9MPhyovB2yclpQFd4cv/p0hOU90mCua5AL1KGi5wD1
c2TtUYreE21NpE7vGnS1ZV+OJZQX8MnWuLGxvzjnaLVV/m5S+Y+AXS7jdow6+/envOH/qoeSK7tu
A2S186hYVUxoSDoJHDagqjWqiZblPJ627rSWXSUWQIdvRuXFdKtIZforCVnSegQP+E9JeY6j4NSu
/OE8aFyqM1TZr0gVWLVeVHFVJXSROUIz/Y1kFF4pi2cCtK5ojobbVzOxfZPDVv3PmxNCGX/zAxY/
JNj/xzYldRBphKf/qMm6OG5w5whIrjsLFraZUs5ykflOd4U28CoX+2J/sLrrjttisCSDka4vhHp1
3w7qp8TEN05kpFTUaZr3jY0MPTTl3cX5kSYi85bhQGv46COkGUKe5CZ61KaHOuqO1Iva/R6lvF1Y
kYAgQDGQYboiIWmwRI9rnT7MXFN8AoQ0ZWq/uB4Lml5FmwjhkMxS7fy3jRhrNxAHP8qffppCVUM7
eU4ijWEudOWTHQU4aeeRJhn0ObG485YVEd3BvI5si6PFnnvcSm+ZCmyu+LJXfb/rWfGaiumXuB7b
F0mZQ2ud+BIuzvombIq52UeZdbJLJ5KC0CKf0Ix37kjjsTNkqNW8ehUu6dg9x3c+cSwlj/XiaX2u
Kpxu8cEPnJifBgjVjn1LSp7yWDtQA5rHmQzKT0AMxgPZZ+w+BsL9dtyJJMFjWpDeVv0cM4Zspo2F
qOyrs6rNRgpbEAst/e9upYo7nTO9xXn2S9WSn9fH1plwf6dQv4x+1iFmf2ds0nqKms0HSBv8qOKO
FXlyiCnL565GwXEMVnWkMAxO39fMHOp3kFRZUEnNNAUC7L9fc8WLg/fCNpa7glFFnWmbJtPXyM3k
Scbwb+lBLBkociVM0TUcI2dkkeIR2bhJbYD10AQ1e7l937q6s0omWRj30z2KyOt5lNY0DGAIvoFk
atUX3K8+V5agq9Qw5RoVPqIWUh1OTrMR0POj/T9fdbgaYCHFG7LqcKt8h56seiITZtd++vqL0Iin
CA8i5CNaqSskfqOF6iwn1JzRoQFuO4G5xMyXUqVHeVbQgpCEo2jHqUWXHSP89uSsNkJKIujl2Gjk
6FIZVUkkJKZJDyMPr3SpuNOArUilYv5KVayFTkCAeytSPN3Eel5DrtxER4LFwm0mb4w/TgwvfApN
MWJ+9UIb5vbwvjGDHxnnIORKFME01QVhlUtIE2nUchBdvPMcnCzoXrf444+LdAe3HGQkIcpxUePl
Xi8rkOQ2FKsTO7SFM5MgrYvAuMy0KAcB7tLPk6b5KtY/ralCMaqytgqkmW8/GQcz2YXRiLTfGTYr
QSNxLVrcK0WTj5I+aF5gWd9Ig1gRqsMVUdyVBbqwhtihlA72ILpwmjMnJYLQz2ktNA+4YukO5Ztd
duGH0/uPyjKEElQIzrbSHmRc6PIfwp9lPgrFL52m6whGBV11pRxAFAgDQLUSpD4stscc4s/0deRm
XVzjLQ5vSV0Z2B1AjIaCXTyG5jpk2vvS/MBr5g0ZprCN6yCIHoMQ+WmEbWqfXUIr/YgUtAuZrlb8
of2wpgWn7JU+JnnAjDDnSARwP/LtZV4websb3bpGw1c2sRRPSbIrpevDgZp2auLJWCkLYWI/HEXa
X1J4Y0wD60sLPRceUKYOhSHG/yuaFSr22aD0RNVUnooqb1CZ3Pf7OPn31lz2ceR9U4J92+ENyxh8
CAOvpkDLHV6pmR2r2SXekek7mu3Ftt0U89Ao4y7Wt6FJPFJ9QuAONzGIIkxKjfyAUxMxXaYKUoX2
IH23gtPd5Csoi3uwjn5w+/LlNw9FBSgXp0mDgj5mHvkqRzA90Z5BdGwNxL3PfsZFLDPU2Iaa980g
6pq160VO+lqL6VQdtwWRnP3zcnmBGQ0Gab2IpK7tB/Boh0Lc6kzXwXTuCyvISjr88+IOPAuhXn+h
nQEV7lBNqxokVwB+S/d0HS8xfr3vs9f/K5k9f1zsnc0azCHNT2tdFW+76Ijhiwv1O0T9OiHc4hJe
kTF05FLPpBajExpv6StEpAQcoQ4a0zZOcU3BStkXI48u3SkOI4NQc6D22/6F8u4zjrIgPl2Lvgx/
/nebgB+o5Rq4cTkgeH0d8KrLiLQOxqb966jBJfWjaml/pQcV5R2IrZwUxMwSNwgq23nWfypa1cAU
NPtMCEVqIIRQSTZMC6JwK7Ou7FQ2MIYwmfxBzWC/Rd8A/5y6+7uCnoBh9kSUt1Zs8eIVuN1JFeF2
bnzvfv77IcQhd3VtTYNadXqlXVU03iOO0jgmpmjkJ06zz4mJmca4ed/jM0U6fESRWXqPfclqgfWj
S11FAwyOYf5r7/HfKp6G1ccPhEKwHyzPFWyauk3xzDV9kU7DLVpnyfTO/+IgxUmk1PowVL7Br7Vm
XROH8H8ntn8TnQ+nbBmp8DZ15d3KJA7aGiCFZToPeSI/1NWFa9iJnZiVwzXG1Pex/oErNDiTDLDE
iSaHATkEmrsTTf+uMeqhgqPdMTAYsC1bcvTHBRMg028+haOdaZlnsLfAoYQjTXQ09J8STmC7eqNd
xO2FOd+zQMfr1WxpqHuyTjGOMhCjDebxxZzsgB8HyM9FhUXYYfOx+p1b0u0JG/Maz0gCBCpGRyca
DpB+8DVpHBjFbHRS89mf/aZPLaIaTCzXrpGWv5z7K5AQq0Pnv6o2yydbBV1upydSF1om9YHxln/Y
Fupd+UBuQaVBcpcKYTjrcpQ3BDhY5tHGU2M2Ezd1GnuVpQRErp2PfLvDIHSWSDaBTSAUY3Q9CbE4
dKnR3QuIS28hs/H+nybX63Onu0SyKMua74wvlllYbvvHuVdgXbnQl4Fw0qAC4GcsoIu30/Qa32ui
iydVk21Ts66bV8DVY85F78Oke2+Ltd6rUtQlh/RCwOv1PRyPWY7Gi9JIhHef4/lcov6soIw7xUNv
GYeIwpecYRhsny91qR4swD7/zaqJxY8gg0BTE5SQYIqNw/cJaOH0kwC33Dinl8odgKWq8HdU7tpZ
GFECVvRAJGMBwOws8/8Ot5RGT3e2SCiMmME8sv1bXfueIoSy6n9sNNzbDv6wg469/ekWVmyOG1oU
WpZHwpFjCc5Fc3d3kdGiu1cYIh+cvOjCCs8i66uSxkYGVVArmnuQjPUaRPQwkLk4O3dhbHIoXx2I
zoMghFGDLidVdfE47rNFfNW/dGkF0bV7AnOELu2QZColEwRsW7E2negKlW1WDhMYHriXbFvaRlex
vzAGwnztCB7GvtIyBPrfgtUL/xA6OfI1aQ6DlsNlvXHZLNq6Ma1YS0bZA5YEOmTRzzClD+AoYLr0
CiTWQxVfau7cERAknw3eQqwdPZmVmJgKQSmtsuqSlaYiUD1o6woHRrbsR0xzXWKD7ZN+sBxVBxUK
31WuiPSb3F6yzsQI3zIgoxWLUmBWCinrUwZcdXgnn5M3LHsgiwAxAbWA2oJrDTstHLdG19CvR8VY
V7POXrJY8rSJOpUZJI1LaYIGzcdN279nxxVjg18/679rRWoINdAln+4zj1167uUOYXL2oeofSn1v
kEWeslzPrbuMV+QduwdKKztUkzFBztPioZj4TnJ8bQQQLRL2KYt1UwH5rSzzQcijp6+0VG10xa3c
DOnbkaLuDqylLutxebPfP4EkdS9d3Vt1T1aP6PJdomGu9afZKHNRXWPbktVUUoCmNH90Q78Fbwx8
FZch4hoDGssaIjC+CFe1Su1N9dp2D1ycQ7Koz7ruHLMb8cVPfbuEWQvP/sleNwI/IKxkmHsKEi0U
gf1wP4vc2a4SEkRo0x0/4NK3G/9j+k+8GItv1nsRIxMKkP6i31XIWtq49n+8qWtUy/aPTb9kkP0Z
484632K8uxQpf9DLZfgoY7bLq7W3COhhFteh0k0CMpkgaNZN4UlyKSJ7dEaNkN8MnM83sSV0rZRI
5qnR84Og/kNvz+ebQgxWHxuVywW6MK9ZvxXaelUCxzdtFzCXSZTIYf0ypafivvUOor+07WFtnTZO
Sm0eTeFc2iV7jR6jocMSuppDVhJlpm1AlNylA8nZSl0QgsuDS+CW5mtHY2HGqE5ZM4sxUGVMSfmt
kFdJF9YrZZGvpzZOB1Z5TDDHwTo0i79qmd/yBP1nMhSU33uaHXaheCKOd12QLdyw/PdIzxoJeWfg
oxGn6oK93MF5bulRTf1zSpO3/3XcvyHorm9GTWchPqyj28/7FA9AR3hHkJ4qS4dD1fz8jPQwJhrl
nynyeLN47f6mZQ/VCVSrNLrqv9ByAG0grtMc3sK9uMTIIqT/EMQRhmK3FExyVJjNLWpD2+102Gxq
AqsIQO9KPDwcrKWbbsoJy0oP91cLwUb/GSpJvexkI9cq2Y2GNtQyslybL4tmW7TrPgfPTok+jMu4
9rgPKm1Va7gkw+DLWEXZTPmNcNWF/hiza+fPb6DtP033EShg5jQGsWUzZlPEWljsTVQTGLOpFk1t
xHtHZ/2VahpoXG4RrtwBWPlrLNu5mTCor0OtBXAjbOd4Ho7owpUEJshlsIakQCwKBw2X24j2ehdX
wXv3WKd5o3yG/mB7e41AIbpbqN4rOnPTwCLOJ2Y/nFMyiw123BeUpB7R4ims1P+Mev74DbtlRKio
EH/Ir6AvKRJ23oiCoHIKh6RC8FfJs1jE1TUoT4ieUm3YpZ2xGOl6F9D6V5Rw2rNIsjJ8GqiV6fbT
Ct4QLn28TQt8nztdRDJsTDKo1JNhXnAEVpyi3finT5K4mBdrObLOFXSX1S2btzY5ewc3Jm47gzym
7gYVNfY+fVCyXzMArSgL6s2k5Q7OQJ9q2rC2WPFlH3yVjUvLvdZ350uEtTVO8KCTUOLDfKsEVajv
5IKPTbaeTjbTWpebX2PQ+p31wM47TQ0PT59gM4EVNJPPbPqDIvGEG64lvPjZNvCkYyX/Nfx5N+CN
UR5DgaiznUdqUnGDjyYL6RKN2Q1AFvjgpDnAyCO0IR1h8b2cCouQCXCaym4vg4hx9lgkht4YPToa
Hu1K9TRAexs4FL+Q7xllt5GSD2+2eqOPqLYEg2C6az7KH4C39LrL10DuVAyLoewHGPbmy4r3GYrc
chXlFXk19k/p8gyD1l7g+z+wjXD83vSfxENn7EMZvJS3sZ1sEffU2OfHGmQwx/atkV1B1PGmOxg0
sqrfCuAxEem3zxs462FhVYT169W+FCarpGeaVDSVmvOx9XixHCaBXfeAwlTvFKN2a/elG7tZwqiO
wRNSlL+PBfhPCGBXJbSFthO9/jLMmtJDN6Dz4jYqiUDaLVPUjdVVe7KgXVaO4TIl3QtLSf1Ocp67
/SWLzOOSJKAjVTOgrS3Vj3zZUpBsCsnRngkjJWTo2E803KSGvTzbnpoyrSiHhzzzP+S334oMDqWZ
H4p1OxL43JXvPrseKFuzd+Kk5HYmJwpgEPHYiGO9eu8qDD27sKS/epKXVXOVdNptantVJo8qgHdA
rrClyIAP+dYKmuYAatc9jX1q8MX21L2GWEnyT35ABeSy69AsT2Iv5RMv/gO+aOUR17kfiL1750Nq
VbtTGSKBVkiwkYsquvqI1dTv1m6w7EytLwd578HoMoOTMZzGHCbuIlF4ySiEQI1rwAOUTsDCXpKa
hZ44hE68bysfankK8qiW+H6rcP1VCWy/JgUSl0XPqH8hApy4ABw/dRMG8tzdnRGKSX8+kXpKlKcE
4x6mOjbXDvTGMhmCS5EvczNQ4hIWG2iPtXn/T5nF/qu4eRIr4jXOtGQ6zs+uR1KPpO9ym2/h7ALU
QiWdMSU97YP+i9zENoGaq11o51I7pKIfXxTxwVerlDbDkb6ahJF0eOv9o7sUmCiTxqxwB/9XtdEV
EKrnv8fJZQOU06va1/zXjuuaaK5LjA+cOhuvcQyY8zUCi9z/chqPM4E0FQdz54vX8miz6kCrHwUE
/uveX/sHX7YclbEVH2BBtJM6OANTtWROsRIhzrmveXUYPULSTARIPyNsNEHHTP8oPW8SMu9cUBWU
VRbpRTW/lXgtKq9lHkE1dObZ37Daun/vPYywHeVvSERVnveqFBXTAHjnyPaaNZqCIWWroIuFxxf4
JN3KxAxrmeWnUyvAGbh7iLmUs2Mu9wT5MOt2uYIwMpQxn+Ev60/FvFpB5MaMnNyWHbcSxFAHaNai
e45aFOKSafSCkwE1cndvomC+09anNYi+hpeRBFvoTQUucsmf5eIWxp+WPRqaBTZxQC2gcNqTLvx+
rfwt8glcHaw2XaF3lMAxhKjyZ7osgHT1rHehtsclDknPxyGnhXDlK8rlm2TTJfg+1f1E5IrwiRT8
BBJnwnmCjj6nYae2cPk5j5HcMoOKESdbtYwkSZsgs9XFTjPqDkiQHgfUBLGVSqkmTC7qSwypYxhM
CaCxLQWxJzcnDeev5E48hZFJqwJGsD1+nsILw6kYOiQkjoa7lqeiUvTQ7e03WI/U23b48uq+fzLV
d5eRK11JLgAR7KmeBiVq1EoiKWMbDzlyVGPDqXcMzw5mMKaaxP4osLzvpZ5YtQ8WAjrE9hoIV//p
unhGIkNvUatv7MDT1FBhkmSMNGQzmY/yyd2OIutOMWNEgZPDS8FMGw3NaGJJN+q70vGwDqzP5dPU
Bx/9Y53NrG1t5MAAcFkcu7eqNw2499arS0eSupD5t56T7O+mtmbBIQQKKPlGhmQEGHtzy4nDEaYd
VVejkRshTmxWeLfGXlolVk/4wbIlvcBkLWOQ8KRXZ8s1gltZKz8kIc/EuKeoQFdMlEFlmmkDM4qY
Y2xT28VZvKgpSrlTOqBsvc1ja5L3GZzEnwlh01wISv43aZyxYRn8DRJwbmk/hE1profhiMK2TvKG
tMFc4fXr1zQtCKsWAMpdN8DBFwPrPwlU22yK35MUcmxvteN0haK/4oYy2LeVghYtUtSdHbecZThm
Y1tmqLYbs0IijclJgwJhOk87FuRcCVG9m4tTK9S+RNM0QzdwuG6i6XQMPFl/ytoJWdXkqLVyyrR9
8Ikf54X6TARdvTx7vW8gaDc9lyL2qJ0WRXn2ZOnhbvweN+PLysn1qjrp9FdOmuIRoYUkPEolGiCa
Ut5n60npaY8D1ze2wLzS+IChVtAz4YKxtHWY8GAq5eol4YHBI+YeL+ve3200E5HUY7jEpVQh0IIC
5ZduOpiikRMRUGqC77cnkf/o+wM4bV1ljP3aUXFcIeGh+sCFsvWirefoGIcSHwsCWvLMYKc68JeA
mpRgmnrGtvArxH8cPGvVSqVK5U+vKltFLoy7kVrkLoCWmVdv86jlAgiociF/uRotq98qQTSpcoal
q0FfD2Q1llF/JjIFLZwkgH/v0nenne93yydEtdSd//SyEw9H2fO5efqe6tggxpto1eYaV01RZ+My
S0zpKknKoSRWMaV5nEGF48V6fgaCKC54SdRjJ0emEWIHK+k2E9vnHXsOukixR9a+NIR7YNs2p+x6
wQ8PgskCSOv2G0vvIizHtGPEyXZd8CJX4RnYHxB7adUbpGfzeTypAoUEMO55Fz7SaG+INLjNvCRl
j9YCzRWQt51Y/yuA0AZ5FDE4WdHT8BeL5x1nubzAQ5kq7AqBOihF4ctTANDC5d7crwijd+rtOrcU
BrFo0v9BC4ueulVieui8k2n/Dpj0Wyv7GvHYefSkR9H6bqw/0ZJvmh4oCFz6nhHIXLCzQFrUq56B
j7nURYeMCUrMdXFN/jVM4ue3cwDS+ExpzHs538LGESNM2od21WnN6Wb4BcRoBeyXF4NPyhS2k8uw
dNdESgARrOvWcJ7XvRBKUBMi3zPRttg8tj1M76iEYyS+1XJGt6fqvRL2UHhgRgVZb+pWX3amA2ut
Tn+KPGYyUy4+AeYktfV1K3h+BGsbFyUEcAD2/aGAvZuae9dKSHnl1FmVRgvQP+KmFNPmDCRJclpr
S77vd6qi2kp4FFgxLKGRH7YSg7b05nZfoOahqRfEHRUvQGi62vdwhTAXRF3SNNocrRUGMZtIPOf7
RYe+PeRt/aapOGyqCWez9Fu2Fpyie8SbFbcf5SLXwZibFlkxnZhpdT4HnwtzcFrhXd24Axfuqp8J
dgwOQg8YprrCQ0HpdScBDCNe8WDO8JUcTTbTroHbg1VpqEU70jzf30ek7HAJiW5Pt9fmhUMoen/B
R3h+IE5pJroF1ZUh8WoN3xtab7Wdn7w1tQA7lOcQP2KY5T8rZn7yXcbB1CWUzPSzMqe0Fu4UwL/m
uJg9tvDrBCPRMsNrSpwQQ7wSIXUWfGx6IaF4ZXcoBoMh19qfilHJoLpukCF3cq62ptw+ZkCFCF3E
GICUL5RYJMGQEpxODatkkC3VwjOcOxQryqlJFw3bqTTJkiPhjOVZW+E2PUSqk0Nv9XidY1Hc8h/T
4pUIGew2mVeR+EOCma/zWbylgN7o1beHZrpyeyeuA3OR9nzu7tmDNdAi6vGlq/ZK0RBJ3xx4fxm7
ipBw2k/vqdEuC3QDhf2mL14xbMSXHcGEADK2sQU12s4NUQAi9JxbuIgSrvrPfgnVrCJsjmfH/fQb
W43xSCZYjU/JtAoua8KLGbxgT0KU6WWmyJZiQmjtg8p0693+HEt5o6xXpj1E5SnoV2Sf0DXgBWi0
FTzr5AuHwVWqCVFCxY7TGRZrYSyBz7snAUwTJclioin8ORYeo1tZitwytuqAw2FlRHbM30NlBRKN
3lQ/zs88kpQJX6fnZVwrwoF2ea0/KNMxgKQCU4ojmxA5hE3qpnU7FYjbNJ9OpWHh7VdcLyT3nmiS
tugD5DpqCcoq8mSUcANezk5lZ3cDA1yD9vmfTjSOPEaxInwz/g45DdrWpbEKeBxoeYP9Ys056r4H
kvWohaOwCS6WIVPNbTGIbL74IJr35Y2owW0YnqIeD6W5A0QkLo25D2r/3SpAw0Hg8GT3Efdm88Nl
IyytMC5FO3qXVSblqhyauJuLSUfiIo3DuxZH7jy9GRW13KUQErV+nY8IWpiecu91pTcJpPaXrr6A
pmTQzdfmRTXHInSElmIE3/SG1lbxNByuEGa/2El+h/hsBUKtIZEZhXX2HD5fI19FC6Ejb099eD5X
+7hRpNufh25UenCsNU0Tbvc7Dv7OIkkx1JMQuY2Drwd5nFqjtXGqbYpbeBA88GCaRrs4TIk3WHAN
fK3wc5LbQLZub/Yn5RQGdHxEPyM836BLljU0WAlO6zL6LDAx0n4JJWsp5XI+aSYIq2T+I4jTdm6Z
9bG9BWhKkO1IotilVZPnnsyfuaWdZbHozqLFl1k2j5C0jra3FgforQGBTBLyDAkcLCHwn0sGbMKy
KPlztwwlrYEmJoS4av1fLVAx4jVrEk8LOpMtEfjcx33aTEYEjxvr7Jgv9Qpd5Dp9/j/bHXDruqZr
t1NknJssK06K9eJvNgEqi3QpA94sHVhHRaLsfepRugZ6GBrRKFuGC3kDg8OHyjSUFuWkE0Faw9GZ
NDXMfjJkas4wq2pLoLBBkTm905zCqafQ8ZLheY2+ueVvjawb1UglnRXFPo5qT23qaBJKhxgmgwhw
DZHBcXNiheD0U1J1mid4lZshZsYUjob0oIwuu7EbUx/Q1myW/n+sfhZ53ghCVxBt6/O8lFpBuIT0
somTRm1uBFEi4qFWBQxRYSTS1pfErQETHImvNCXA2tlPgLvCiDRhuiKfKz8w2i9NFkn2matj+HLf
o2SUUeMX27id+TvffoeMrJA6gXEi+J5zi0WjsPJByejaXSPapktrEwyguUpw5aw7yOwP9hHkcdzl
ecOmu9WQDX4R6eFs91rNYwPOptmLsUTCpca+b2maHL/ngVMv+nU7cohwqCw/6+4jDFbYzR33VmAo
yNemhWRcsGE9r+PYU14jd7B1t6aje6U51a4AVMHhFdje4hio7Y+4BUMCbeAATtNnFxdun/wYNX/X
U20VBupTglcthnK0Zpxan8GYITpIvgnFwPJ14cs0olMHZVLeckdnBwB9QtHMoceEuRn91NQRrSTO
KsaMm35k2zI1Z7fJ5hy5vVo//TkB8mNAYQCFFaywOAo6/c8MD6+Vyrgtt24aIGqOQeU5F8aYG0pt
do+qcVrSWRWxD44GM4Bjbofbwnho1hniDpwchyTc3vfbLPGpIzlsqTIgjoAOpbfmuW2KfrgZlqdl
xK6DkVvunZl8YgSozeBU5xsr4/CXFFT9k4Cbiu3apiZR4S685DByxYdO1UPFcuJtJ1Jcb2Lz5KW8
8BmHKDQGkGRK5xvYfC5DVZJZLwjkcnNQv02IUNKXEeDLOoginaoXjEeZ3IzIscBhp7ZUbQsBKCXa
w3JKVHwEXXXIzdxTgO++CWC7KuI/HrmUovA+LjPGrlOP8nUrpojwi6fSlJfNm/APO1uqgX0PBf63
uxibelCNBturGnCmluPyyTqd2U0o0MtPJqWn8CpvOnJLk60YoNmdiQOlG/nKAyQJyIOn9SG7SCI9
+5Iu5hom2upyhjFFY1supHtnJDNeCtDuSlpYJcgF3Lfib6MWd9xdwmNrN1Ql3cFaMtaaIQxg2dZU
+dwQ9Cta79KBYR2o+K/0biho9XJF5MFqEeHl1KWkihG5v3lg01o3tAkjI4Rj86xG9u1vtOAsZMgI
h8TzmpFnuVe34q4Gkb3gk7zWXQNzk/xt7mye0Wp72ZmFYIQbFnuYps3Whh90H+V6ypwjy/nGYlLV
8eCbVu1gw74L1Hqj6nMNmAWXWyE32yRwq8ThhbDdAbQ942NdJ/+CadH5bjU5PiT+1Jsd/RTwO7XK
bs1EvS7vEKkjsydvBxtU8LehNGdaXixaWHjtzoUoG4F65EJYCeMCjyLQrwsxKy995/klUKMhRPqV
d/l9jFXy7illIesE053cZ2/6Uc7J+ZCoZTizN9qeiN0eRSjZ0NpPJjhu9ICVYViCtMqEZHp/bbDq
Z1jr8ZEDfUwQ7KdBVx5oJPdz7AeMvZlMX7Kpc7rIRisB5DPvXrlpaQjVfnq5NdqYyAPK0fv0yDim
LO3eh7OcSb4yhoX90muQORndKjFqEB6HF+Zb/Rg/TepFhZv0GdhwpMNg3Pr7JPRS05mkLG7agexY
hSn+JYMio0nZit9xqXlNmYw3KR69POzZkH57XVTjrDMouhZY+D8wF67Y7wqk2In2kea3SWsFQA09
vGAJTtbyP0hEvZCNk0swzRM7UNUwQGfVWaq4Ba5LaivQSTFnXrCn0Xu2OIecVVDFi+C3+xwrBJl/
iOup1twxDshOCAfrwIVdR25jgliW/hv7UBV+W6b75o2mHID2qI8wHTyX9RX0/CJMcj4Rf53M/9RT
wWq70wz1E/J14s/fiPQEuDIMt2l6Kttt4AChQ8k/NBGZLdffEnJCdIoAiFiLujSz8hya5jlQWp/j
aUNysGCp/X87I5L2o7N1RXkKe3Y3DHanU+rHouSQLhh29WxrS8D/qf37adufbdySBEe6lOAsds1I
PKnTfyBvhMywDQ6L5eSWmDCdaXbEnRneSDJNPArE4UhCowlA6CqHbolSTVF4vP22XeRBpvZekqWJ
s27D17uszJOMuVg6rSncAKhOwiOMNalzXpMDTSU7c7evJT4D+nBaaMFtp1jjjIy6Momn5pnuMUuL
V7KtUqqSfyrfC3CguTZ/qBtoydyyXNIgg7Jue9hLn5yKmrxL+12y/xhYmcFB61/KhYJGB6yCyXka
jVP+/GnB1xe6irCVSjAzKlpqeiWnG6ZfAONQ4FnFJ46AK97sgFXslh+vN5X/5l9NMB+7lMSSYq4B
Tw0i+5AD9hdzLBmPfQ4sUKfHKgYxAgCMBryqc4zI8+k/x8okyYz6sDssTK+FXVDD1bWEvcJ58cJn
NHq9Zf9vwQfS0w42Z5FkncwqIupuiXbH0SspBl+RwEi1fZCpyIda1iJ0ElQofceGQQBy8jQbdeVQ
wuz2OxnU7MD5cmRguonDDvIwTAgtJLoJLLf4tdOoaL6AKZv1NpSyX/EVz1AT2dzee5xTKLLXallP
JUQXDn7YZRTughT5M7GeHnMIGyF0cz7sfn/rq1OX/+DoX4Lo9I/OiEcWs0PrAEIu7Gr2WY3HARnj
tKnRjFOc4LBKr8QF5aPAIZOrZB+PDLC3xUKRDq4pTL7UCMTnDaBgD8mLmMRKIS/Amw9aKMRhF6h2
9dlYsc2XmcTJ/gSOZ6p0peMvqmYNxPv5C8laP8q7G8NrYkKqNmiqK47xlQHXfySMK6j3vG5r1wMa
ejiE2S+NH/cd6YWxf25OFR1RVTqSmKMIK+pUkraldEowFN7PrI04YoOjrT/1wY2pm6dqXh4zONE0
cDm9PwixzW4J2qtpQsoasktJFKMV3x7Z2ydSpefypuae0GaTRdxyyG4KzTNJmsMwcU7bwkcc2CFD
xdVdIK3KiG83JZpmJJjrEum1RfOtqMv8pvEKjKF20GYLyJwEYlJH8yzwMj2yl+ryASXtvDitZV65
XayZXV++wkswT9W5DjeR8OMPOsYSBtbFKzrZjCiOer1qfPGpqacaRxMTTd0OEUG+iriyzMHwDigp
XtkscXKriHe2xWml+/G1WM0P9xVRg4aGCH58el+XQz/1XWKL+Igh24+YChOrwvs1tmTm+/SIS9sP
vk6unDZGZgHAJSsl8f3ONkKRdH7HvK1MlfZ1Yo/28fSkHkQ3b3TYzJwvsnYWRq5a3lQU4F+fvHrS
JlLAWp9hoMbXA3IM3C3MY4fEROftGnXHle7dOZjvWMioHrDx9K3dOe5mvblcLrvAx5NFZocOCciO
wu0U1zIXpltJZxmaNz/sygw/5ZsMs9A4gYsZi5lpDPQoO9vIHjXzHYAe2ApRztKjm+zbRTEK91uD
TEM7jBRuKLSc3m0jJH76uPEH2v1zVREGv+BbnoaL/LgG6TUzVKBcdjimiZ2dXX0vi4uKfNO7xqL/
DIZ1pNlC32nFWa52YKw7pj9PikppcPpHg15rAUigbOYVqlArQGcSghCKNHylLFnTSv9yvUWJYpum
OpSHngn8Ks6qAeXzzkavCd1xQuYJGGYmSziD2erQwQWgpPYJRk7wt4kT+xQF5TmkCcYjKeaxwEzC
kpVvM+Rw+08qt1pZWTmr63brnZ+hvd2nfDrliNxZaoeIhWNAKKstan3AebNP+iUI+rAYRrpuwKV6
3OGeQFVItGPWaU7aR49s56SisvAfCLTph/W2Lwi18TXMeVaEVt4x1f43c1zW++uUiePFzQXt5KvE
fmjSzR2fw2wFHkVIPCYUXddjSf8hpTgQ2FfLz7A8JhL9dpBULlV5QfGRH7M+sdYarCjkEE8MKAxh
vd72922I0Mz3pCLmatrx5424IA3DKhzWzunBw534Qph4Qwd77IA+0ju0oCgjZdj7Z3Z+K/LVBX23
GXybFd5pE3HB1NyzEc+l/+XofJQ6lGqjG0i0xp6VcDM11ya1ukpkktVUbWLDVubBfXX1FZRiswvQ
mryoFOdNveOpKShivD0f9tHHqsahCI4oCesxIlPlg/fqgIiU3IIdiCzn/0y9f7mBDfQ36jgiv0OS
jEMN0p5Wkug84+zDAHndZURBkLOFNEvZ/ZbwAQ4fDsdBCBFlpynsiA7YlLzTeIJQfLtAA15kctVG
1kHbw6gLGhWu65SztePAwKaHd/RFUhv4oPbGWAQppfIeZeH4dqfDEnRIESlcmaJjukWDINPCCJR/
P6gizfKhrm1+UqEj7bweFZlV2qChz/0uhe1sc9b1vEuT0nhN0Siqe8oyA0MONa4RhhPVfUN70Qgh
n9e9OzssHzC1QSA+ItLgA5GbPuvtun4v+i8ZrDDX9g6ZFAQd6NTqQpYSgQbXyiXR7+GEZjFdxqem
fDKNAAZ9HIVii9wJw/2qFLl90xvGY3JJX2PSzCBfx0ZXBHk0l1unHcdmTMyjbFYUkTIygPukm5eD
vWcr1NYGgEZQr49Fd6RxsaUFR27uDOQ23Il7uBsWNUb7N41CMScCT9y4wsaEnCO5t0muRIgJFYTk
Yn72aPff0/Xs8UDqUAzfUsANsRMEoOxw/qkO4gTsUYETl4Z5kQlNxrRtmqiYQZf5fKLu228Ufe/5
ybGZbarw7ohk1HDbTLP1Ciuf3ou0Q2XkMgCQpCGTctKndii3Da4imEGuwrQn/cLVNCxtnN9CMmmr
/YdT1KiEq+3UZtSxRblv8ye6v2GKNzeOccSXEbtx6SLmBtXKKVKjqq8f6lCev2lwVWYZLnG3gUPa
zLgBs6DH0Di3RwqsF/KomQTYvTtkjsWcPin8nUhhi21y3rqxo1YYwklu4C402NAo3gQDTCy4Up+p
EVXQOCtRehLIRP1JxvKPAMXxm/ThDX3TVxvh2E+giFiIto15UzwlSkeb1Kvq6Y++8mrgsoI5Gio9
CPAFfH4zOg7YaQYk/J4DqmzUAFAZlpWTuNL+wa6xMSL9sAoYvPAdhR+ASHoqclZ36FByyeKVRy5R
OvLI9Lu6D6FCEXGEYYULXP8Uvp2BFZbsQEaWdwYFRUTJaIIi0Qd4xd3vUFhh1kWv7RAlSWu0rAjo
QBQOzJEZt6DrvxHJ0zHntCji95qG4gfbmkBNFyZ5nFI3994DJFmViPJrM1lEn+Aj/f0mox30MJYG
1lr5TxTZhjpKuOPA1nhos4MHEzBS4tzWXXpuJlkBHuujz2OLI4j/QEPaVOjA91hgo66cSAVc82ri
QdalJAhmCyqsPQxuUiNOeDk4pqAEPC+eVKrFLQCEcFLtLyKdTu1JC6+jIhlzBsFU1pLODsxQe6rg
ibiuI8nw0f0R+6zLmKL8dSzCwsacFbDT+AfIIoJaHLEeaaMBZChHP65Sq+71PpgXu4HmN7Ocdt65
nMXjU4JlKV9IwY84mTc1GHA/fx2fk3OOD/snBk6cI5qZxfkHeC/wu4tkRkJ3OxLTD+pCcjFa2boa
YhC7mwtoaSuNbalkChp7l3WrIqFMr2RJYcaxoJkqQMR5XEqC/g0o8JhM9VHiwnNTTLa6pLa+B4WG
wGBWGIIadI6rco+cyY5XY+TEkttDltb1I9dhDTZeJUQA0/UyGR71168j1IOgZJuiUkknDTggimbM
6yVLfEl3SFQYB9nWS5GbrC/OMJjRSU44Wn984L8YWEoh7kgvac55/VisCj+BpYIkIpyeO5yuRToZ
oy11gc5Fq/M+YvRBwoldhWhIKyD9vVmQRyqLsEIppjq3gIXebTTN+WsBRj3domfVf87v0VEmtpMs
pj64onwxKZFmcZ3lOKn4ujsuqDmAfEjvdSsXy6SukSYgo+YLNSbDwEoU5fbBPcbPuGkkljS4QfXP
4Q55KLqfkfxjO9vWnIWnCu99lrHYOk9Wgh0RDNiNYV9TOIgpwsycp+qIwn7NuYu4TyLYdIfPF35X
uRkKPmquh4rb1Es0KJytXlrjK0NmqXISHo/f72bKq7v9vdLbnGhrW0oEPKPpwqVSY/LsrUnvAw3L
jpyMTmdnWI1TBKLwUdU1P1+sTC2Y64aiyKxqnSZnetVO47xqmpRiqAwfj0Kd+DYmdX8Zl4GzHv1s
ZORW05Rd7pTeOmLGDOVLREGM6ZR47I2befiDTvJfmRqrqtPDBX9E/Ao17s5sTBZToOSi4RuN+ZvY
TgGTGR4+MVzYfOmJuebpVqLVTFZAh0qiyXl9h+2TsUbQ8YnI1CranK9YocYkGOD2yE8tFssGE+IM
EeI+ofpetrFLxx+kjFBp0CaBfnBPKHx5VSRjPYgzIruBJMVgL5WXMS7L3aeRKo6z0tR+pi4UAuqP
yf8q1KlD0SpIb9jOXQthY9DaiH2h5CR5jRcEcjHLPsieUI1QvwFS4wkWxB6v5veLAnXx/yjAbuGo
xVDQIsrRQ74tskqzpmDhSPHgQOI0oBKSCWjUrPTY12BwTOHs8BpsmmyJqK8uGGn6ggDiidaD0luX
+r9tCXV5hnZ+9PL/vmMdYzBVOVISuo5vBLHdwj2DmaabBSKNqWHEXtp3jouEk7GFnY/1JjwXDMp6
H5Fk7I0kQgstpDVr601ieDW/+gIq8NyPS9Ws7SV7+8aYOJ3kFsMwUYNPwyX6xZsVIpGiGlZFT8Qt
ovbsjiZ0M94QmAskVUKN1ctObzp0ZqRFTIIAhi4dpR1lM9mO6B8+CKi6EaK4zXi5VuLJAiON5E+k
1WeL1uMnsxO8Ibm7Cg5gYKXo52YeACoB3Nc/p91YbT/+et7XZBdELsg6InsrlW0GOLA8OayX1Q2F
Hqo+lH4h6LDyURUCTOxiJ6wVyHM2Gq5a/j4/mdgPjCBu3+n+l2sABnZKyxv7VdqrwgsdZmdyL2T0
eZ90cfLjDQTPytUnC/UnPwHxcm7+ehsI8b88ysgwkK1VloYcwberUKJ1dmzg8zwrRZ9EHuU4KMw3
4KRk+ZD4Uyy/U+wqingIS35AzPOBLz49GnV5R4+XtZmox1G+9VFVj9nHhBW3mIc1cNFwjOLzP/9r
UTW0nexvG1PlmD9bwXw+hVXdLPxAyzu8H9OiVh/+n2tz83SN1GSKhAarNQjyOwCke4larmGRiuT/
oc1OGuxkrUv+7KzdBmuKEcxNmy4ASCDxxNfIkSN8CBeSha4UYyYREjk8oAvta8UJOPWATbEFH2Xm
xduAgznOAKKvjxGtxKuVJjwrY0Sd+RVGk8BHQTok+s2G3YFNJqe41+3Zky/iygBsFQnHpizHxhlA
z+smVLQllNtTi3FTkWxSLzP2W8yyEJv0r1I8Ng+ye425m3xi/4sAVvxfG8/OEaeZUoReVXAmoGk0
4P6ILIduu13d2MZuNO/A1/VHqsUWUmh1JmHVpXbX0r/JRvIUqD1eKrNazWCnyok9AGBSPwJmtED5
GBvNYnhFwwjbFGuGnMqN0l7MrEK0fOudjhttz4+0iSnpzJXtVrkr7/+Dqf/kHvSb6thQPTGeaBfh
39KEgRe9gBSgbCLw0JtC7QbwJ2EZU3+ybxtYOm0QU9kAC/w/u1HJ8GAHj5kBl+dos3Fx0vlz8mZ8
NPHNLj42+9rSgsNZEqCpsrfsDfjyeEInHttM8l9yo4qhsrwOlX3rdjVCSVoXWC4WpUkx1w0gmRGp
Qh0NRnwY3xnOGDyq2Ka9mz75ECJlySLpj5/Ql4uMxUKXIS26/CYZXy5vjlo+ilM8lXL9B+3gOExU
9p2hifK1Y5MUuJtQMvyIMDlj0tTDbsxyFPC1OQGc4XijXkJFyk9CWm8o//LOP0Bgep2D45RjWbq9
koL4/T9i4wgigGON42EWJuzhoEqkUN8D76kAbu++33nGwVzDyw5Q+f6B4IMkuFZeMTyY7fPFvD81
DfIZydGciw0CReb/UxWFGbZMPJExSpFQjdYMyfKbSapIwCdmEnrNgMLGCGH5v9c6tdu/88XNwv+B
5RIeMzTqcBtvT0uWQds+8rhzdkw1db/8KbjaVCWHgVe/E7/M2zJaXJ+pgSGHn/d7zgLk6vgTDQdT
WUfZIxMIAIxMgimC7QIibw6nx17eyUsCLrgIQ+5qPXm/iNprnTzjD+G5AOuM++k9iUQag5ltbUkW
pDcusC0jQgGuf36ouPn0P06D0StLy/iXWoQedWur2bmkDUL8tQohIBkS9TAjopn7rW9qZVV+l6uW
3qypHhj2Y5YWF0R4wqm7vDSCjnyZsdzMobCY9oH52AHUOXnNpuUDQ44JhdH27MVIu0Yk8k0t6o+t
p7jM6Eq2deyY0deJAsgUBMwQ9p1m5sxO/rhnBYA8B75e5S5bjrFef8OfC02uKaFDY6AIrKH28I/u
f/q5Tcd0V7rLvguEW2zkEnVY1FmVyi2YDeLbqM6ZPB9ohJgb2w8ddw1vXR40c8C9bYumtxEOeSxZ
/RmMshkeuqcuUJd5M9GVtjXraenxuJSxFrwvLHwQlCawiBbQrWUaR8p10RDsYhMsSCDm0cexFf3z
ppzE25M7nmVqu1L41gbvMtNdxkDGG5HYL3wYZ6qmjw/k53o15Peg1JaEASfTnSK526JyIu44TCH+
WK24w8FbDSaKM4EKh81AbmzaRM9oSsJv2ag//5CQCYsAKf8aCcLeD32xseZj1C2Jz+aqxyTT3E7a
YgHZRNxSelsP7v4wXJVKeB/i4E7maPKtXiX+UOprpimJbCkVIltApeCRrwrAYRufhtgSV2JD2csI
DKGv64X9zzKDL4pplez2ZfMrkvW2My8X8Bkgsi/EHTwm25MvuHqWw3VPb3dCOcbjQqeDU8n56V1G
PFmB/lLjatvS8jXFYZ9Jx223WtXmxXQu9ivJeKHMaPJhucHhP7nhcaOgIo3RW7eAHkO8r0kTAts/
IAzXORqL6SAnL4DBkiswGvk388SQwJ16E1XsRs/pjYlbVcJxUPz19sHMSsUhcpwUrmw7Xi+L9/8c
6+hpEbveG/Mchgmsl+CLZGci2XotARvKJtpMIMIZgLD79srTHFJI6Y+595Q1pa6p5L+xmHlMsXJi
ABlpjTTIc2JpBKTmJcdXovZRfUi8mzQpZG3mgSc85HpcdkF098eguZERD/jHrlQavougRJVAlWPC
bjr4ogNqV2v44mVc3IaBCRl7l50qqklVlittjrp3HmKssntg01MfGfIrNmcGdZf2a3pG0a0GviQF
1glHn6xTlzVh7NTJdkwJFm9X08tzsZleqdk1OKsF9dpj2hdZbAOwpazmHtlgYHH8hQ/xTsI+XJgk
86cGsihNADU2RKxRbVrY8J1tAoXM5Lc1GWKDfBeaf9VBm09x6vmKL/gerixRztOoVRJjxle1vVU8
i9jQOt9iizQSDYxRzuzS9IbywFskp9xIS88SqR/hjCeAD22FuLfMFevygdPhMOwfs46oNYTwbNdm
4hceVmqeQ9yx9bP1kAgTko7EJHzbvxR19NwPNKmjTdOgTco+44H7f6FX5te3VHlzAzqev30dRNay
SNsOtQTRnINz8ZRJSsGJn7nkOKzFgwTdGdr4lUdKJXtL909D1M+LKzU6//I/7K8YuW28E4K1ODeS
VpAeyuaaueKX+HTuxXFGLed5bMiVZ3rtUTa/85dyri7CAsNxnfWBr3Tnmpa+YY4yep7am2m5e9Vz
GnDLMkwptRs6lf5I7N704GJR+/cySdaySaTgWmr/AoCFzKequN5aVk/8UaXVO8l8S8Y19HdlPLZK
2YCu5vf3xHTr2LZ+6oAE3TN8UsWevUYcFCxHVAJm021E6kaKx/xRaQdHE80bQiDY9rc4/a4M9Ugy
m6tmBPRngrGMNE1eMsZV2Z6ArqfBLh77q2PaSTFzBckjub6iijPtz0BBUKOyMN6j6a5Qx0BOPMg4
kSZ27ovJ/Cfv+yGVWhNOktGGHbQmwMjDGolgvpIjUgXcp63JX12+ZUtilPmN7Oa44twXIsMZbMC4
SqKau4yqXVxdXIJVUKEsJKYyTmXuHs1Tg8TSBjX7Kc73jOl37x4JinbCXkd9S+PtAaYtEQT1bIDi
aGBLnUSzZI0A6tY2EuJ8FYeSokw2plUA2ZtkboXReBCEnsGSEXW3lHgBZw8kFYYla8Bz8IpyqSIz
OOmDBpBbSxwsJW/Ty9axIM0t13ZSqTtBDA6LELnPpLyTCkD82gwR2jpsDjHQnMDkBra34twQA4uM
XTc0lG4QcFQ/zSNdqpHwk7nJIDueDbmCfILmucaUX6SxXPWBu4Wu5yh2Qfm7PyNgnEj/+lSklJxb
akDSnk+DYM7NMXe1YRjssHBthk7gMaXuJMbapiPPWvjl7TBAPnl/8okW8f1tC4VhfoeYWWQJ+Sjc
RvCF4MG4Att1xIP79pc32zycGXJpXogML1C/c1/sENto9JVE0A7ny4PpC/f0la2lVyxKLxlHUfZI
7NtCFjXSDglUeYe8i3eEBQUPdUnleBZLvtaTE9WQVoEQ22ydmdvVsvO549fdA/6zdVu2n2G/vey8
+JqC8O3zzwenynTQASyhU6YCrMdrCHhKoHYF82j8C27cR9zuQQNuG0TerTeU3FeZouc4hQ/BoZQQ
4Ig52CDbAQHbqipzmZ97pv3YuyzekGuczk0gLP4MTVko7MdL+vzzCWpt/eu0UTlOPYnG5XhOcZ+y
9ihFP4a3r1NrEhW8ZrS8ZQMGrc5lNG9Bfe3RUFnFm8GUscsr668BFGurE+199qz2z65GNIjiOJcq
cmEP6lBentc9lMuWQJbzuEldo7U3cb1DSY5H01Df/FyGcbbHUnjwlHO8JE0a1zlE2hJofI4i1UsQ
qKl1SpuhUUMOJI9A2aak0hX0JX8eKoN0sVLWATi+/prBY6IefVR4AKqxqsGuazMRCHFWK1ckoSrg
VE89oNwykU5V2c1fsSF1lTUWtMoOWTrPh9mzw9yppZRQGjzV//h0gTmi4LrgHae9wA48sWvFQx51
I9e/zXN3FNgSedEpVOHKpbe2pSKYB5wEKyTmlE5ivU9YAf3TzVrzmRAPV9DU4NT/uQA6Mq+mPfHk
OFmmVIM9ndXdGHD6uYuqGVtdMmNf8muQOQcpn5mXMUoUFzeNwPg2FIKlzZaUzcZ0p7uersXSFetr
iVpvmBv02aIZyGYq1U6nYBOqrWS0+ltwcDA3z+AtaaNDCUhJ7vrWXX8FK+MC7W2CoBlcYVRn3OcX
arZpStwKXCg96yeZU8kuTaSVlK4rMYS0Ezlbr5ab4tq169/9mDl54AJLS9W0RIzAv/crhJ4uPOY3
ROsZTKr2aocj5Mky5T1qQrWK3hkTSlucOu99xNYUByl70bA7bw33qxM8+npnS1+iJ8/+4nrU+mES
3J+MKN1rnBzMs0kdc1zdfblDMx1VHeNjLkmERpy9NNA0LpqbdlKpV2rdBMb8lA5aAy8WbrVtGqnk
N7YZdewo9FaaOPEinhTXsS2afZlDubOmcDi3m90Ar0UlxZ2izssUszjXk6eKCCuMaIuX56kHZA6/
bBhKRxhv6rDzVylbvgnrKFyhn/IkvAN6uKWXe83JiGyHDt6Qz+CevRL+nYBQAdmreOEj8o9NZ7Sh
JnsC83XMc+G5jpStqUSH66TIY8r9RLoO030SHDW/tFYvsEOb7ENEzzhl/Uc+qKUIjOS8crq08Rm3
Co/kI7ZgdBP0xY1LUqt++m3pvEcLGjWpSRVwdiGr0Nl5pV1beieC/to2deyTlhpwdMAU8B82MTSm
AZxk+nxnZUBeyqM95lIFGHBHg0ZPtziUMTncACK0krqUN17Y40GD2y32JdXnVEHeoXx4AUoeMXV7
jPLfQPTdXF1dlFOUim5yWgpYFrpGnyvoaQXNthJSswaY2sRLRf8ZHdeSZZZ+zFrvh68gOg/D6Ipc
ScvJoNt8IodNZjdoAI89MrgiwTUt7gpRNgXFtV+mNnEz6KeNvqaBt8G1w7kcIaj+Iz02zi/ErNXA
9sZfrTyiu5yP/05UyCFSzukIgYzupz3IFfXhufBX6VGG5U/cK0yhUYEpbtPxVa3o/zIeZMsXPDdx
8x4P+yxw/FpPeuyb+yfkE9h4F90ZHHZ9tYmgEMvJKvE3w/N3cgVKNzo4t5DbOxwFVm+mOFULfWNi
Eqq8NoKkhfM5HQgNZv2I+klxktlxEMQrXcRBvY6PULV9scT9QczbPn5Vvzn4fnabJatvCRJThS0k
lRm7OwB8JDSAoFiaMkqCU92uiMupTYjVhjODc+Cc01WfPsnDETrfk+o0wA7Lwjykgtb9qk5/QoMA
Un8N2SRyj/GXfzow2N6zzrf9OI8p+W65zbJOSs8VkJm7cY/1oMFfN5r5UM+Ln089wr5SOi9cCWZs
dH3xQd3Z91S/quj08oqCA14F2Uzwj6Be1Jph6xqJOkptqlOZNBBdq1i3fSO2cnnUsRe8Kn4xdaIe
Bi0I26SsOdU7eMRD3Sqvx++uwN6b6cDLrozlOaItSyLTrsoZ66kU10B/RsAK3vIwdJEQ5zTQhOFn
YlIVPybmfwSxB0GMn8Wj9aNXbtQwwF8SKjZWcmOwHqd4PL4AonWkvRxhQiUJCq1bqtH6xO0Rq7K9
MqElIFV8AZgNwxZbdgYitFa0tQLVsm395QKq/20aYm/2cJUkIMdbt9vwJ7lpUsS1NgQlGeUp/ymd
DXkSTxzfPSIyUZFeT+hBCHOKt1RKyCgwRct9J8VSVzo05bY9w8VufoKFR+XE7XrtcFLikQcR/6UM
U8r7MaWXIUv9BkQX87yEpJajrMJ/3XnHsezOtnarWgq5W9mm5FKutkkC33cOqZD71p+e11QZksm9
4Dpjre5qYui6wLZATDTbmY3CEQd/J8J8dl3JF6quxzbqipSAShprjDtXqguvToFf0Zg7JtE6h1k7
sP1IqIqFT9rClEm/83ZBDb9bDQPhI2scTody0TyCSysuEDFH27lfxqq3bogs1a+gb5FgeOEBRnGh
AU+3F2An7c7UBwVS95l5MFBFapqTIkYR6mzNc5CG/Af11WmZUT7SqnUHpKdu0u8rwyCZJmRw77YY
Z64MTwNzK2N3PQp4MfzeuJv4tr24WZQTshT68NKZqehnFBF232+m9fG+p3KclJzNhbIBikzojBHq
+eaH3n0Px674oM8uYTSTBrAHxrp+xKh44hnmj+eLasRuWeP4sUjCtKsW3Y9KbEdh0zcHoqpTQGiB
010z+jhlAT7URpdF2zql4KYEr0nX4UtHUnGUSG3NnDXmLIf4wVmcowLwD0ZA0S+xijDI4wCQ32sW
LevDmV7l6oLaqpKXOMwB+EOVyeIAt69AzB1a2CAKk+43TnExxBBFfh0zH9TpQioJUHV+UCk4swhB
WZzDA9JMMme3umFu6ZSnQCzDaQzx2PEc4iyBVOIRaep+4e4RQQ11qsUguD9nlzPJFf+25ricSRy7
emwVJr+sbwVHLn4X90ZP7RCpNThl/yL2mI3/JhHFq6lpwphBvjNfmsqP37En0MnPuj4CFZLpMKnR
SCiF996jDrDYFmjjjrvOl+3cFgKZh/bcu32NfHj6anAnx7zxpJlO8K8eXEXVYs9Ls/AbiRxJiiGf
VcJAn6BGB6Od8cZRzsfZnjK//tTMSOzN9Frlw8vGnUuY+d5GuU4jKQ279ndxW2vy5Z0M2iQ4IbOq
71/KkMJMi+N7WNUKij4zebS2DsDokVPDCRRBtdap5KiglTgIQOBO5TUfvb6blaDuhtT8HvSp2RPy
+TM1kEmhlglRomkEflm+1dNUuO4yrI7650udD1RhJ807CXGKYgJ10PEPQBIfpD9gwN7MmVaGQvGq
E7z2lpaLyJwLfaPFIIBRAqc13XNFsMoHgs5xpAZ2buMn475DwHdQpA9qwdRhCUaR6ui5jDo8/Onn
BT8GzC+3ZQ4Cyp3XehlbGWIsTKrYvHiutyUVxGMnbPznHF4XhgX9wg+itB48515yXfdlP1UTRLr+
O9PmKqgSfy2Zqd0EZYLDIF8MD65iNn/GFR26vWWUdVji0BxM7TzH2ZlgyCqryn4R7GNPRWZRg+oY
WBrzX3jrNWtIOrcruXW49882pLbizTTySnH7hxHs6P8Q2g669Nd3akbo24mFo1HTEmDYdxO8fX4Z
i+1/Fkp8BWxjsaPoJh9STC0pSJmXdn+00mDJI/z003EiL6vLVmcipgbih68kAIpHM8XbuLF/92hr
z5xU0cswz7fJHrJDfsdsBRaEH7YI1OXJ82cbJqutZyXkXwGiFexEQjC2pYarEVPYCW0ByxxjNqnH
Xdg+2DR45MJrpQ/Lp0hdTclFuoYLmr/lzdkATVu/rlqUQ/EELjva5BAYzaJTHnn2cZmnICpUY/oC
5l3BtoYG8MqZRhSHLgNe/k1YeucE4ADc7uqozlDTIO9gsOttM30O5GnIiHBr9i9PSRhc3WxFbPmW
EY65mTHAx/+YuUl+pW+Nzsg8sAA7ftyqywuCPTwemk8cZPnA8uti7fdMie1/8c2rAxY93j+/k+06
PaLsvDV5vkrKpq/MQ6XglRVuBsUyn++Q4zqXEMaKdOsvteraX/Yz5cn8Fl2EXhMp+owhyMSrZ48+
85hBDtGJdhxg54uuWPwJ9ozw9BfrN7jt+3aB7LW0t1nROnsCHdlDkhIytVRvkcjNa09YqhXcFQLk
rWFlsVxHDJ89luho/67jBjoy5+ZZAhgUyWX5oDYcJPexkWh5/08xtSz64ocRiKUzVeZNawyP8jB2
UajT0eEnp27iwwD7Mq7K95EN4DU/XXJv17IUUjzILN4AvZONNJtCw5x93ap8AhH5DtRaIKDSW5QL
dyRnE5187YCdzp/QMj2dnotJTv21SM522KotGgXE01htjOp/0bLwZsme7/neZcjcxe3s97Q9cXiO
szWZDM5ApCWkAxcQ8cqToj5OhyI6erDDOYOglyKdpBqNlZQCzS64Bt2ICaw5MtdQPGabkhF1hEDE
vjccf1ikxSAeWwLBkKIOYYBdFDyyaIEnuXogYv7sbuuhC2MrzFn0T6MfTnyOrnjTmzMfpNaw+z/t
UtpHd+fP4Z0iCB2Y/NuEcQ31nD0uRMx9rM/XzKQY2M0KO7aOUdbeWe9QH9AI9BAW9OH0memojgFA
AsJtLD2f1gMyF0Y3/kfki3S4WgUcbgZxfibRtafZ03GsK450CIYsY4qDIsv+cYj+3qscsHLsG1oc
RIzLd2RfjqhPGTCVi1ytVLeUV44pCbMcUwXnvP35EBKanrIRSQyMWsLGurAm1WmO9QLklp9qApiA
K+At22gQ8oT7see7PtGWtgDQzgemLPEOz46P/EOGUXigD22Rl8+SXCeIu9QQZ2Adiwuh+x8ivIHl
VuM2b5XPUtq5xcwIqW0cHvNKg6T9+ugoEMIOBRtyoRbaHy5crqz5ZLT86PW1I+idl43LPZB3c2Wm
6pL3csMj722FV44NzD382KuKrX3hZGWU3zz/qbqSZw6uPJN5qBsrWaYHklRl5taxliM1ighsf0dJ
VnNMIySpGfguUYS8y4GKw58TMv7w8DYHpcuDm0FSq49+mfaenrvfe+D5MQRHploQeKdBW7vTmZ1+
5XW6ThcTOeHoNEaWvSAm2fP3rox1E2+RzKnPf9nfZrCdo1ONA2W1iErpafnLhMXLfdRBVQbn5E0S
M2HRKsdFrQehbj/tmwiN7g+a2CW8eP5sxzKvNoVU1JqwqM7HKnIwVNtp9wVgq08DCo+FgtfnMm84
AFkKmojXrTvQc2koMtR32o/d1uMzWytxj/5d1ttwB3710yDrQgHPquWOmETKirFalR8yNjmFBQfM
AO2DH6wS139RlRTcHTTgaKY+xLIrcMf+rqyEEWxQq0lsyKBHyv5dcmHnDX9Srmlxir3ZRRge5gL9
sW9GDuS1/EStPOthApuHiJNJi+4CUXeANc10W3/k9senDXqGk1a+e5SDJjN7uCnzoi6NT7knUDQM
RcseK63WP8Za2rXZZK3+aLBO2NMUw+0QXKWuXebc/nWldWOQ7XanoeU8Ii0u+jsf25ErUpDBu1gt
oYLHdVdKC11Ts5i6IjgfWfzE/O3wQPbAJa8QJpsEHHxfZE9W7j5od71uMc2Vv4B62RbnMHNqGmWj
RyU8ZqB2x+dVgLXlo83q/AaSIb1QaisBVlfTjIuwqVGYyCZj+TosNid0lMYatuOSTn2x1tUx2kZb
CIsMpc2sx3vxEejTinKVS9SyCx9KVOI6p3hvc+q4NwEPydLv5uG89h/nVC+2wZsMp9Iy9AHmScqA
Nd6bqNodeDLszVpsQe+mDuD+qnTLUJjr2dlW7HMo4o4zJGRrfCtDQV6F0dEF6xn9xBYceS5MlkJO
FSlQLU1t6kkGqX4YU+N0KdaQaFSBVCU+g2r/gQff3pZYi6sSi5sSjVMFIFQZrOTtxguKQkdDHhkB
4PPhHCBgzaYJ0+VC5he3hXMampWP6hi1inPTECIGrP+uOrAa4TmzpjdJ1La9CIc3sSjNxUnwyR3q
s3mxOXulwU++Ev0iHaKrgaE/Nd/KHlGAubyjPX+HREp2TeM58NcMdJoQoFSpkhjkGIWOgDgAEcJr
FlzHNPmnn6ElNDkvKhme145TtXAGZ2UB36wiD0CDPQaGN/MtZ4SPZsXRwzg9BMgPeezWL+PivtJP
Sbb2pvbAvBQcRyUwzOsWK1wQz6KQnaFpPhv7BnJyZgq+aTT+edBCOxuOnKDTJNJjJcbtASwLZLf4
7ONisWy1VX18lCKXBVELjMwyLTg3UKQ4ZCeyxdiPWce2lAXvnN3a8jeVJk8ETTym6Vdw29ruv7Ii
RmtWrFplo8cyQRh97ynRHW40VENxq2uQXkXq8zH1jYAFebb1cANylayI5INtkR3d5jaNck8wqXAV
0eor2nQ9BgRpG1uRmAMf+CcCubm0fsL0J+nCTvtgH+nXddm1QWS0LVI80dU26cOL+A2puHtvIWMb
IUIHyCv1Xh4XB4/SaG5qrgfZQRGrFiw1rB2NAJpt2WH7jyyBQL46M4hiL+iI51KQiLX6YJ7tIrhb
4lhK3sj9pQX5nycX0FAoqx/5wAeoszgeZN6NHKstin6OwBWI8Hen5n7iFmYCw3mbvPLxEatqIXjh
sj9H43O0iuNBM4KBejocVIS0SNE4aTwffWoEoHzhIWrWo5VYyzkAH8mj1VUbNnadI8jd2S3ok/2i
B1kycg1H6FukUVR4rZM34GIIplRI4sLwd7H4xowcUdW40FoQekpxTGEHun8p3xg3C1LzSLdg8w1T
AngMaGKvWcSzFmgBaFAhjEGNxFzhioG/aQB47aj+J0YxQWf0kTFJLTAgoVXp1ZA9XUOSmV6VZC+Y
Q/76Wdjb8YBM4w9aPYx8sQJTSnZ/ZRfUveSJcFfmaM3o/nr5fputqehAUgpnOdvVAkJIk+44MjeQ
vudP6EY3tUvc84+DZR0J+nUFfHPqtOssyMNE2aO4+/R3wXTLLDBEJndLYwhkwRSGugnmYth0+u1d
zv2UygCQvvq6GdXDiUrZhayTLfNYjIY2QMlHnRUQwW2dIhlucyzk0VAHrGP/wgvw2X9XEmkGp6Li
ZVV+8w7guGZr28wGChP8jecB4KQF6ejT/kU4WQgzBSKCW4tsUwwAvB+RywnmerBqMIc/EbCh70MN
YfJFIG3dsszFStfBA7cy3px8zgVG+Et4dZNma5S51LRk76p1K3ki/r9CRBSErPUaH7S1adFUi+Pk
AiQoALz+qW24nGkvQ96iw405SFSUZNERhfJInhPP+3+VvqriifCLkahTBonULl5y8/qSDMwWUIF9
MeIz/7EtvkPqbz9aHgo6yhLQQTncQTKeFO9HgmoOateMtHHATodsE1s1RDca9kagIV/JwIG22oUK
EQYIuvGFrn4LJOTRE8QZzNzW0thsDw7QLEnuA9Uyrc0GKxhksWglbekvAbJLN2zxifUTX1WQ45IP
V4/JdO93cTTdtpxveo0C0xVOoLo1LTWJGx0hi8fstLj/kWRouEr5mSYUkEo5/AKv4fVe6tU+oxFp
SUp82N61ZehGxhtvI5CdM4J0Z3AODLCpyyjg2twJzNaZF9niAQPSjAbn+qlPfTQTfwe8jKKRgLne
kGgu/W3Cc5817NzxExBfrA11fBNxKo0oH1fw5aCJHVVX/1KFXCklylR6bavcyNR3owGjugnjw49m
Y70o4vM8WEPw30fQfGTNe5v8wGuosEMBMW6YzUoFEoSSvKsMIvmJQlb95dTxSZ5NkALysV+Mfvbs
ApcLrYvZsMepGL8AGOtBQ4jOWZthRvpEfifBeSBsWanXzosHX8mxx8OXxFdHHoC4EXXzxeVRu7M+
eWx2c6nfCOB+m8gzl0fZcxyTXQB98xPH7H+s6IPCQnRe8/4wFAo2D7lIZ3Ov4NeBQl9D2ioPOg4q
9uKdNXDkl4TG5I3LKTEnoq4jILUg5ICY5pNUHzpMoaLMWpR/hdhE7dbyXYx5WigSsiZByrY6Vffz
C5rjtHL2ixPTuhSojYERMTeODmCInODMcBgm6GRhN6xzA/vQGUaO2jA+jW2fts07IhGMBklahSl2
NSwMS9kgXdgj3EN6IAVvPy19bRQa2kRL9WhqH5jTuFNZW85orxfnSu/exlOvgnW6k7ceRCkyzkCl
LhdZW0DV6cVzbM2FavzPbMC6tnXNto09jW0aYsvDBYkLMQZyA5SqASFcZ6vHfP0rAzeAnLiZ6mdi
PTlN0biQUfuIIIJZbatYoLl8R0ejFBLM8pdkaEtNyxsetBM/8aS359f0PrBF0pquVVGPGaFQQKJi
vY1mNtmMHv3r1lP/CS7yVRRbjRpmtNwmarmvU7MZx3JNSH8MIllUTs1IfXI9fI/sfNCTGykNm7ll
tjwUGrateQD3jbRKopCfqjkw4xpMjvgk6sds1XlAsIz2NzFxRoLnj12Fh9dexpn0ruuiZBrr58q5
ywQua+lXYIiwbINMCcgwfzW0VON2kmTwOIYCoMtlBzEsabAACvOkzCD8K30q1UkemPOGb3iRGQU3
eOFb0n3w5gi5//LqspaF5OedsD+/2phmvRqkl03H9HYDAFF4v9BlOqmdg17UoSprfUUzEzu28Wka
0CvtDDLdMESO44v/c4arxCEpGgrwp4xX/eBtO7mEaB/hSN4Nk+s1kIVKnLstT1HCJd88Sige9L41
O7xh0Uy1v1VbK9jPZjwvMwcWFFMDpNryew/y/P1GoUZUtfep15VCtPAe/wlcJOEtVD6rwdp4Y/0z
HIBNaDGEDZ/B7BedPjO/pQPEp0qstX6HypbLDJ72b2V/RhZc/3mFRtEn7EWqGxylQLHXkh1X8sA9
4h2dWcvh3e+d9/BngP4eulvqsClL8J/lt8vab2bdWDBUNsbW5Cnt9laBFuk2jcMYg7N46swyJ520
MQfAdkWERd+R8PUmq/mfDimQd35HnFNasXgSFd/VbYSxTaQrSU+gU4/+MmumxguIq4FfF8fRjj7u
CNjvHRILVsuyjYfrLZoR22G6G1fUTvDOkhDyN5TYUdh68RPtxFF1UNTnYIc/R08nr2L1RC7BtpeE
6ahGrvQG+y4R9bYMR8lBVlDig/aBTFjDsVLNXgvSCGZJfpOYtgs0FZ+nGBXTC1dPLMIALf6xlkph
2zY4+Lnde6Y/RO59DLz4UOJiJomxjtpMkbuLKqOON7SvTkYZ5/rpCDMZpHfItNf670fM3Ii/ylBF
YeSM1uoRX1/ZO6Rq+egb4ya4ejPexXuA1/O97yn+IlSy9psk2naTnB6QiC4yxL5snKAcIYdyDqD3
u0rWusLmxtOT3E1qn6bei5FPWDFyaa6hccgRHq6Y9vpYmbJKS4P0M1qVROm/JMs7qOLs8hmLiPOw
hlAvR83mLGzQPqLmQmF0IN71DcMJASWpLSr4FRc8u7NcFDS4q++zJMqa+6EN6dKDOTokaKrMO0R3
0wNhUVh/00H22/aBNbGTndHqNGwHQo3HkNds1ehrS1X/EthjkyAAvhRDIVB8szaoD2Kmp4g/5sBR
cr10p+2iwZWZgZvcZzZK2IhTIsS+KAQml3zX/54v42QaCoQyMLDFtoiGdQxY/xh4aWrUeiadqe2v
ztpTgLf/MAoo9lIBDQ2/IuXc9jGJDNXLCwrIrVHTvlBaKCQP2KMRoICuQE2migqJsGa+wa9o7k3u
uDRQ74OwHE5aAtm5B20NEEAif3nHD1pA1K3vDPN0zTBBUVw1jWx1AVckLG70x8/uYRW769LmrQTs
DWjKcUr/d1j1qT9tcfdkJrUJFl4u9lk+6snoFNSDONGI1fdtTnhFoP7y1uw9Y0cBg0z8NfFuOzL9
iGXtVoy6x36GpT3Jkix13h/v9opQ67+E468vZ5/vfkdLAIWkscsdW761D8V10T2NLxavOfNx470D
AvM+0YdPCrnrm21VouSLulRDLwhDzV6v9AODqhSgVRg7MUNruw9rQqmUaH6eZzzFUlNfTVBPhc5B
0qy+OgA2VrqoIaMvS3oE7weoPyDMqDy+l6x0mc+7JfwbdxdMJHwg767mnec9GR7HnLAP4OGWDn2z
MPf+mEFs/62IYXImzdTXOkmy/jh9OCQZqa9qaEk7u73ccQtywanWMwhOSYjuq4lZT71GB2O5n5Ar
l8yW+F0Z3gpmKZw79vIgwHP40TTRRn6V34Zdkq4EeVdPdHOin1rLwRMjMKWMowxEPuCZyqZ6Msj6
rViBIg38sRFG/gLOejODZj6qkweG9v3o4tPwwHUuRcTu/t3vXdtp1ubk24Dyzx83hjQlPofm3GL0
sn7/QfKxnwJqIk2BVxeFNdkRRT5lsmkFpzWIsy58fg5irLerbw9kpRiitH/fScgqHGqYmk9cm3Zm
IvHkmPgECjkvxPXMGMasv04IynchhcVamlYV0QDY4bnED0xzXHsjvTtfJSlaZxE1fPKvAAqzL2rV
Rf9+Hja0bq0+tLPK0zk9O+L5AhoNOIco6oWCnIjAPkaGlJetQLs7c4ewgMVnkIuA32fhn0hWiq8r
0MFW0XLxdoZjKQcx5z8+7XyEDorrA/8XYNUvk4a8p4URHH+ZmO1BQAznQoEO3/7S9+vM+mlSNMXT
yUU1F4oHjBSRzEc39bu0YCquG9bekWFmhrGugg4N/hHKO77pla9pkwYP0Cb/q3KKbjWk5QFRi0mI
7S5whSTbEdRHiWKPhsvfLwTORyt0bmLWM3hp8Jw3ivvN2iEcnfXN1dxTfOqD5N6HremZd0brvBqw
Ue922c0l4iEkiMQKpkZ33+662ZmQFqypoqeHGySSEdwcUK+V7shrwmR61Dmr5rkbSklhwoQbGyHu
ygrrfsiWaG0Wn1Bab24t7a9Kipa8OIzXKdpe2eHWza8irLjFOWVJvc6A1CdFOXdsmn88GTKaMGV+
uwllkeXx/zeXtsMOnb5++xatUX6TabZg6iBHmH1NYeypw2OxjXTiCa5Vs1cCUSu6o40KbwASQ39D
PK/c8ZWQOlPumxnWTJxnUBnEFZHYqdNADmhmsrHyjKNZ9WVK8KXtm8nymk0HCVu58LFYsrdU8U1+
3kADHupgIjMDxbLdtTarjw2KEiqn22V1N0rNdCOmKE2q/n8RLBTM0Y3U+rNGF6l6MPhGdh9J08wn
dCydHczmhqmu7RSbyd3rKZtRQwVh5rLeo9FcHagObJEQTtH28V4p5Z3E7YlfyW+MZKATyC6T/MnE
m3XmjbizulQZOB07N+kZGB0PrbKzj1P12TIDkyiRFzETBimgI3xWpc+PXScomGtnyd2XxjHgCEfL
mBqXw+ws4MXqND0XeoAN0dYJSMMgwwd1XKFyRkTBXlEjRNB95n9DbLbI0eV8aAbKFSECD+dsUXXy
ZvbtKhZcJBYFpVQ8viXUXXXIrdrQzsVakzdUZhYahpelbaLJRbh67yOXD/cTCFko3IZ+v2X1bF9Q
RXu5dePHzc9S3uAvBEI5zQdzr30x3xD5nqHOOzUcHdOcDoMBbyGLck2aMkNlkwJ0dJ6U8R5IO97p
NR6Mnzfu06BQstiTKdP4x3h9C7HbDsfMMqvLcVJxCG/ZlLdsOhAoJ+0HljCTXSQQooS91yNXXbqz
+CaLLmwmPzEeOOeEVmRn8ZNbxsi8kfd0XzvYQz+Jnc9W4kKHtFb+DD54SS8JLLSRFx+iHtLX88n6
XiqyKa+RX05jmu+wchqcabfvDOGvImNm+TVnTEU9UxOmVpAR2O7JHKWWR5nPrNrYGqfZQyHJ0lTm
3f9y+W3VUO5sQv08+I/uj8GfcoWp7QDPJJLPAdTB5vMX/+Jl7C+vpRriPfmC6Q/IhHdTFS5PSjeP
uw4PQu0O2sdr9Ey4irddmfzFNbO8/bIHi4xoaQ7anIhwN7IaBNhlx4eDlt1bu5lfjWvQo3VlUXBa
uKlNXpMGFB+rXY2INRdT71N43III3CV8eoiA+z9z2tnJ8+FyIr7MMsL0V43pJRlm1yUC52j7fSG7
T2ANJhtkCK570an54cQWTwb+q2JMxLbTtP4N7hmoEDPrpwOLAJIfvbT5OkHEUggXFriXoyyv2XuZ
HgzJcJu93RIyjN3BJYKd/Q/YIqSW2PVyODBBXKCo6D5BKSpBYt/sYyBVjfUiHMpjTOHGy7KGzuxu
rOSsEDYQMJ/PwY4d1igIRMwa6FiUAVJbkgyVekPp0gCBGKn0W7iYaTso0xqIq3qEqNCSGa/cgzqJ
FxgnWmy7LTvWc1QynMZdmGMUx9k+B2DB5W0epWJJFpHBB5xmdFqtQ5iBmz+Yb2F6pewIemjfFUe7
0lGY+18Jto2/lXD2pgNkaB87XqLP32RGX2Mx6OmAp0rDth31wPH9zQ4GZK20i1/J7AQ1dheYJEnM
I5MLeg91bQL0IOCCUPlHriWXEH+o1E1pRcO63NgGnh/v1upyXcu+CMF0pGb8FAT+R2xuqkdtS7Me
TVCWf3iMwqe7Jo81PfSPZ8lRsn64vz5AqGmqB7IEiuQQmuWl3jrWp0yBi4RZ3kvQmjQ9erJE17Bw
ynJV1FkewB4wvpzEq88DAfpXFF5FFFWJmRd610k8RInqJ0ku6ej6gVM2i6tWIb3M74H334nFC2XU
hewRktgFI7AUIRDynbCLZF9FqZVOkwMm+bVkz+UdkVOUumkBuh9HTLton8W9pkHL0XeP6Fkq1K1O
AXkOKheQb3BQOd71JrF1qC8AAJFer6ypb3EuBz/4tQ0vl1/9tEtUHgzoKLa8L27cP2BFd5/7yIvc
j4JqYtqsmf4nRV7JRAvisN6LOfKcRtsUvYdg3gQajMqMqymtG1PVH2YAPGbAEJYUC7E339hw17V9
8zwNjcvEf0bpmenZw2bnW0xBhbe/Hu5yx6asdFDkNFBUQcSI2Az5hDObUXAkq5PSThoBWDx76UJG
QXVOoBl/IocKyBWZPj0Tqys8sVKx596G20z0BBrz52Tew1uD8QE8EDQlmPiLYrzdwj5Kv9tlQHys
TM6qbc3kN+YebRFrA41dhVy03QOLeNmiCRjhjXJiCOaNq/2V7DRUXbUzPalRe/s56p3fTKtSFauQ
NggFD3Gelk6wAOL9D/JJZ6swRKZkYzNVzjJ1IopLsdbbzOopreYyTkmSMXIFt/I8EdyfA1DgI8FD
i62tiZvKj/+44fkGfZz//JyjSEtD6krDx8canExGhspJx5PWxEZGkH8FKotUHQEgIrwzNU5QgXaz
7ZmkJ9yCmplqGGHRPUGwW+/cSOcMu7pRkF5oH0KUY2kMI+sPxGIKs96DK0K9rKFv+snMO1KrHAuo
PMfzjExGokLTqfVR821FiAj3Cw53Mg5JmfHiNrBBKarLGs3HAUnnybHP1KB7TplBBBBLqrFaOKGJ
if1mYZOOVB07ULMqnf3YQS48ISTPnTNeMTSZuGTfkR3IC/crJhAN0uzr2TYKTxwhQB+HDrMEwmwb
N81nmD5tND0HGgGw+eCYqkrjcnLLiZ0L/V+jlbpaawRtMaBIUp9IQharpRPzkIe76+75W5EX4at/
NWfDDtuxMxzxX/ndtT+s11MG75NoB4ZBRaMvYhBczmtrojRAr7gWZu3u7eaEJGhbB3ce58wiuD4z
Y1nu58tSxg9HjBWl96H+M6mDhyMnotP7VaGQkuMDg1PhCqxypHz8wWpluIrEl5AIv5mBk30caO7m
63WsY5VelzDFz+SeUdrJ7GAYFK0ytd6tq5L2kCXkAWWzeWSDLnaIMcH05jTJrvPRGlhWiFR9Lk9X
GTh7L+QFPjlkneaJ7jljkvN//z7fxTuXXidP1vkOi3JNuPiZzDqu9T2Wy4vNyESgBjked6ZSjUXz
edrbjxhF3PXYXzq+1JEOBgBFbBhcUzD37YsfIrno4rxQUN6JusCrFIs+Q7AOSjaly0n68x7NzBA4
gvylzpPpqdB+sVosIhOo1A351jP9CNwUbj+JhV1GA0K+ZCn/4gJDBz3sNej8ji6kYE9ZDVuElBZ5
264qw9HAjHZXcNiNDA+mCbMNGOkGK4DdT4Fs3cs0zXw9O8wCQ6TWh7vdXv8X8P2zl44FrQCmKfnT
IwVxEzKOKJa7z93Ubr6fI/9CoQoZ8Yj5Tak2485GBIvDIM8nwAETKr5zhAzYe18cEMEFdFNrezkJ
AeYIyweNVRuwNLUAXuhQm+zds1Ez3uusTx+f9t/WOriUWVBa0/RFoMfeVV46YEAacAvYQcYtIyfN
FJduhO6Y74LB/GXikIoJl76HYaphnOCcfYIc8afgx4bzUM1DwZ2BhubBPrL6Y+iOG9ETzdsEQ8S8
dtf+6MWQm5unLxb8sGlBrNBN72yLVrlQccNwbj4BIPiQw8WjrqgOqeTpiGRirsHGkcFaW400GgRL
zC/xdYQznPGJC6fxhctq8G5/8AfZlc4gKXxefyKZrAJ7NvKcUF60omRi9e8+n+fmsbsdgtCKOfnd
jJgwzbKefbRoAo3VMBTzDljoAHVv1BKsa9Fg6UO3SyCWoKj77VhO1NlhfgzSbE9wTCYLzQ07uvjN
KGc5C11BKAB4OUnKI3fAz2TzY9LgA4txi5rorRT5W2Htn0x3MNR0P73IcQ2JwiE46v1tfBn5Uxlw
YkQY+az2VsznZbSLXXDDqcjWwP2J7wxr/8oe8XbLpWAq7GuI2kqFThisgmi5F6NUJsgFfqvDHK5a
yQSlG6Zms61aVSuM5DDYKAqdL94o4urYurvfE9Mf0Edgoo8JycR3yn8kNOUGvcghXR9tUh7ZZvam
ckKyqBdw/nJcckhFwfyirPfRi+Bb++h4yyxTAKiE/NXOvDHZQi5GlHPyIdBg/p4to04OdDDf+gTG
7+AeHo4/aIT4opueuN5qxLYIrjGrf9Oh41ixZOAtemedMqaxv0JImTv/EZmbGJc0K4cc3OsC9hPP
6j8Vh1HSpjanX6ZgEQvKOF4Wky5+tfCTTGS4bIU2DIZzvQ9d1bHnXdo9gLWNrj767lNA7JB5KnWa
fON8FNF2ikFO7CBPo6JBkuU7NuiXT06yv9xg+qTpHfBacPtei1A4dZzhwC9+327BolQcikPmCxqT
kf7y7wJ8dJVOH3ttrp2rTxFVsZiFR5sWQmCNm2XgzXz+ao3ax0jQeGLV5Ubgbk4T19JgAREcJw/+
AyC4Kbl2DCabW8hWFTDBSJADkf58ZeNejho2pbZy5AjMi2VLs3Z0LF2PFekYQuWHBoOMcoNTBUFV
YGKvkYUB0WXN7/ECj7siqOjeNtIkCwV2vPrIjcDib5iVvQeeKVGX1w4aOS8080gVojY8aJiqvOc3
6MGEQiqZqNfWL2LSZjYr5lhvsykxvTGmFwAwkd4a1DhOjwxGuGoU5G5vkZ21VTj7i1vW+wNBo+w6
O1RoRpskeQ/C+guqRu2OY1haMmSXK6h3+fU806VRbUV29WK+Iezl31sU+bp8fT25d7y1ePY4J00S
PwwTUjJ3Xjpxs7HzXe50kgcQQTezGMOcMQYT3K8WtxIpoOIwM/P4RITA9AUwMmk2fhX/aehy/URu
7LkgllrQBb9hFO5rTsJVZ0eBiPmFAWMZfE0Cf8nLt0KT8XKyEvymKhDurVXoze/KwoSI83I7uJvT
KqqEddjpfisw5khPT2sqg1BChBiRa4D8Isg+bTjwFpX30WWE5WmbMT0rKuCqu/oSIW2oSO6xPQMY
9Q7fBaIeT1x8BP3Q6CRbRsiSDtcAifl3mr+hGGaKTeoT/3fyVbcWhwjOHNH6SF2fliZqj/xD1dxQ
DvrwlmZKvxRa4N4NBmXCFEAeiG9yQ79iZjR3Rybfu+etVCmImSJHmqfIqZ0P1C4hTyVefeWKeC4x
PwUZRJlhi9HVvPqPwCEXFJv0PHwYnsIofzdoucRgZNyEwW7IWGfimPCJfWBYcjDkQn6OZYcOp5Xu
Ce1GJOxoVrQwFxr+qTm8l+RnQo2as0fGp7hKjS9yF6nImvuRMmdtti87XcLCm+/rsusjyr1hnHx/
tTKji9pTIETSJD2dGq95b2Ld+nF18m+5q8jtBIz/tJj4jPS8cD4SQfLlSUEVaiV+i5YXrwLFTKwe
cM+mkzuGkrJZduPRIEcgoKr5gI9SbfZAy6f/kBTdTRaclnD2qUtwm1iD7+Dm3tb+y1X2sjPLFsDN
2ePI197hFMDt0YmCwxz8tfYkaLRTwWZNgkH2gzlG6aT7GkrkGYEpKwsspkjaARsQbAV1etsQVN0W
NL5rqmqeQqMUDGYx1bCt5+IAUo8RYirEKb22zVuUa+4QlPBNgBh4zW7VIHEsearqBJVzX2pmOzHv
6XAoabF/WT4/atynbVPi+5S1WwEHcVQCCDcbHVhRlItMJGt6/V6X0MSBMO33MeitToqvNej/qN4+
qthhfDdpvSI8Dx/i/kJ4faOnHjF8Wxcl8WDx7tVnjstNpUZ+Tat42JnW9j09ks+qAFsy1NZc6b+P
Fd+f0DMFAuNld6TAqI7ctyfsbWCJaDJrs1m3qKRTofl6MLgCN5m8uG3140s+vQbJCExJlOJfVaW9
n+nsVZZNPk+1jmnLG4EqWpJ9Td49/aYkwOnhFIYVXFgnLf4G6WdKV82RvfbboKUQKIfYsFJxU69J
Td74jG3iGDzjyF6LHxdgjTzl6WsT8OBT/ztti1yjDSXusxSoU04ARqx4kpuHMZVdIyOJvXcBrpyT
lLrBTnHk7IFufZmnsQhCcQPHnnkahH4hspHDJu1PJ0a5WDH4MWxeKfSC28Lsnrwyf16OGxORHJo2
1+6Wfu3B96iwX4RncWmPjDQ4QgmLD4CElnrbns5YIcX1xEPFhFtKZcTDX6NqH4RUQRI5Yx6liDPT
cWCGBE3PZNLCH70SiqM5+Z3kfcpLef3/d+Y//50uOozjggLMbXAWBEuWm1xtvPolPCIRCNPwVze8
CWycBC2Vq9KOYSpWu2V2EuubkPlku6w0Cxmd0V/jKXHPFdNwDE88kRJ5jM6ne0tkL0Mw3oviaGK8
/cbrm09UzncYcIb/6lhLNZmd/n27dwoNArVCB/CqrxQEO6H/XQJo5w6z0RrsFiHuPaC7ZH5/fVNE
Q0sheUF7MndPEIoBGBCRQoy6hxmfgBlND/VRvMAVpv2gHUQv+aWiIKSCaNLoAIgQuGCHZtR9l3lY
gP/9yDK733ZMaMuhc65SCtDtZiqUlpCNpc1W6+uz5IMe8IV7cQGXrRy6s0PcFCDRlF4a+KQqmEBD
o6o5yAr5hlcO4XkGe+e+dtWOeajDFD8HoDM/BDfJEUtnINkqeo1XDijscj7ZjGVYmh7xEB2vUV6d
Ru4NlzWEG1FrE1b9ZmxJ9omJnqPtf2ZtTBpR2crZyTT8/CM8FQTz6cKukhtojevkUVmZlGgcar9K
V7N3fwFXcZtruhIlMF4hI3j7uk6VBlNiE+JSGP8nGpnZI5gj+5PuZsL+ORnjOqD2tdyAUb61VZzI
t4BMEo8R5eucOcVyzBmZjBkvUtprImH+auBeEb+PDNLeJavdkbDbeE0goxNG/DEU7zyzWiS4+mZm
FXDU2M88NVZ+UAtQCVMF9eJmY7+ES2LoT9oN7h3OQaO3aWwW+b0ttQio3jUR/Pa/frCJyszEB9hW
IoHSIKHy3+8eblOPAjPA3EseB8OMEgihzZg/u6wsszUkvKqbUvlRm0HzEvzko4E/ta+vW0KL61UP
6THrElc6/GTbmXf/0GInSozAoukhs4Yn6o2U9afw9v7DY0OAqLgfPO1HVkJaFP7aRX/SRVdQvEVo
XGAIHzwhqAWwQqvPFE1gfKLJ2qSLAegv2WUR1wpB2gUJ03RIwcH4BAOeOX26p0KtsIA5x3h9tmQw
/745sWqve7FkMEM9l8jY0BwAr6hbGf+TFcz8/gjjE0SxslbL0zxEC8FiD3zG+K4JP7cyYkS7Zzt1
Y42YZU8EaNU8iN1GlY3A3L4xSGJG0tQhBL4DI8i5bnwqxCsmW0tmviHYv0oiH0UDdCvVVp44IfvV
swL+q+JlSc54/tPlwSfEeJ1lzyDcU9YzL2HAnb9Ckk0u0518u9qYX65oLMKqmLPZ7QXZW1rxdazK
OJJBaAOJuORqQgKlIJqQJ27QuCH2zAChg02w7T0K8oAKRcGRVartkcN+7nipLR00VV9jdmJi6mFh
CtevLaqQ4qg1zB4iz5IQRAd3lDgwwdErviiyInhgAXN09wrmekWxi1zFHv6unmtBdL8Nvw8q3pSx
1ZE97UJrSYHVXQjugL9V+xg03F6KMZhJMIMpKWtC85avz3r5rem92l5w2AzeqyqVQLA5VP8it8ht
SiaUJACzpjJ9NaCdWr4E3dRSl5HAUkFd3oJ3Uhf/Pzvwu3cDsfs86QyL3VkCkLH0xo+tECrbZtqJ
y3pXYkFh7n/vJEWS5VcfGHO4JlmheYRbcMUNM+CtZjRyRNPphD23FRtfqDf0wZsk+IEQvjcGUKd1
S3CngjpDgG8g+9YhZ57vVS+eSLIQx1L+iJWkDzVnnBxJqmDW3zwEAklnPIoAuy+pppKyMFvE76PC
0ylpUJp87quaoK/i5v90pqQsadj0qojaWWghfytS1vcI5A6ptoLWptzBgeWV1oUZKqgyJUeS17rG
mrCiyQKRc/7AgU3cJydaESpmZ9pcYmtbR7JocCLrHNO4MKMFgDtrj8qzpOMQfY2aMatq0i6zwdQE
XcU8qLYR/iM20BUB6XgF0CcO1eNMAoHQbpaOH2YcVKdqVYsLvQgBvkVoMXH/KduuVyi6KeN+XFRF
96zmMl52vE+ecnbqRKUCluHG56bOhejpWLlOCiPzG7KT82pOdjDMjN7Csg5saKtCXvqYqDPHna21
T1sKSf0Ias66qWc0zhLEsF01LpNj3UwgoYM9ICzIzix/jDgh7jmsQIpqfu2BnSZKk6uezHNqkUlp
gzLLs+Z9yLp5OCWhZDdmKwwDWISd4nEP8ibYmN28dfNBYGHamPIiDDKYuA0Z/YeID5Ci1eyxtG1G
aK5JT3yYgczVYcpWexiR+EhBvZ10Uq4I/aetYyfsDFe4MUZUVOs+rh6WxvW7srwpi/m0vADyysBM
wh9+zYa9s+mRZ4uy0UN+N2q2PXTHXbvBmAIhSVApTQ+5wKF/shTqgWzazhutLnaLjTIqVH94fwVU
z9K6s9E5RfUyXj1Q4eSMWsINy7l6QzZma3/g06KZWrU9CFnU6MC7oP0Kod3t5yFrSeasb3/84Lmg
lGjnvY8bg8DgiLetTtiBWsvDmxj80caeoemP4KFZOjM5g/H0WgP2XVy2ZawAYyUzKIBCD9z1Sr5p
OPOMcF4FFrebXgOA/9hsn0i/RfNZJ9bHyZeILTShfZzU+Qwo2DLDLXOI5nSh+R2JKgez4w1ht9rL
XjbUoF8v/clBvr0VLKp2no81lXQjoJXc9qq6MZ3TNJu7AIOsluvmmNzf7oHmh7yVQ1IlkAPOcTod
sP83h+34qa1p+9RsdTox5NFbWycNvVbrgM2IXdZmp8TggDcYokJRJZ9y3z6QBgsmwpHd4J3m4Q6B
mgDVuoyZnfadEVgoDZobCvpW4wSgbTeBLM3TF7DDxyz42kVuNYpLZBLQ8o9SZWVotTg4XqeJxtwr
FDtWrmY38h3aKtO/ZoBLBAn0MuEQ7Bvqs7vq9ZBVKPusfTYwuods5PePlGzJ6LrRgKclHjCeGJ/j
isz2TS6uBxZoHIRIlopXY6/jDPMayBVygNT3RaeP3EBF+goSXBsa/ZfnaqqZrZ3ZgV8omgL3ZTIv
hKL6Uph2KuFI0HDa93FfMJ4tg8w4BzXkBxWKM4wpux2tqE+jQFGnnWUlTGaCB372EAeU/GhkUyIv
PHlnUPhSbYJw1f+btm4na//MRUiRwDplMT7egK+kGwro3GHHe/EuUPNociV3vswPQzj9WWhPq25j
lvIEh051iCBorgSGSDEOg6v8AbvRrtuidVXJkooKrAmOYrYq+neQ4INC3c3vcyO7laxEge23jx/Q
6CR+i72Ax0iwEmjz93M7q5/6EpIgARTPgJa4qeVPakb7IFrUSSbDhH5qDLLIPiTpcjmX2HPWwptn
g2lpZGc6oqyj9jYpDW9viTtfwf0JtVXvRwV2u8gc8cguG0ivkcERmHwY8R19wetFPQbpVrd7yk+E
HrpBPq55hYhuHtKk8VA7YMnLwfRNQW5JxLGsGCvYmhXRwx/jnIqLI4mMsPWeNdq4kzRppo3IXMc9
JNsoanMePAjMTZz4spJvtv1EQ3E2NYsuhxTnFJ88t5llCHYagzesQT4PiqhjdcjdQyTRL48Oo1Wa
z6UH+VVqhy0LpMb+qOpc/i4DcWPTUbNcubchbkPtCJEFZnNeVz+Qxb+OGC31jrBMC/ZiV/RpP9es
DNu91C2zjFJNGGyhK1aMzINyoV7rw+04RUcLmfSTKKCw8zurFYrne+pOP5ZX7xQJ9bfsiR5+mjZ2
FrYkx8ohdFcykcqwr802YAwVhw0cY08Kak3W7c/8YX6zRtcF6AaqG7tI3MXaGsZ5qvdY6WU4qzW6
MVH2BgKIknwjjGMQmPYV3ngwpRs8oM+D7OV+4EPq//wVtOzNqkNMGRPO8+dBLLdtmt0vheoL32SO
7ng1H7wtVnyWhw7jqH64DAHCO8pgizQqKF5/oeX+Gmskrpie4epsKcviPNmb58qcuGj288iQqiKc
qacVbEIUTski8vSbzjIAlFpsTtAo+9yR84wVwyL3xUuEhtQOy05I4Tx4e5VV2TTOfXdYLsM4cMy+
qWEH3YGStyIwM9MgU2SS0GlGXaUo79a2oQZy6FUFH+ee6wC19Pu5j05ksGME59S+AP+F/TN0bwen
GVoFHMtxHgoutm0/M6/mDrpFe86YeTQNK6JFgSt9dIcWNA8JyIXDhTnnqPz10u1+oia+6b5SCXgr
wEIosdItJfSNA0IvSGpw68V9dqWLZfFEYVxO8tJPdzCMCUliBrl0D8x2xo8j+FfUVwgMc4KkBgl7
XSSztUQhHdSC5H3x0+0umGxlofFoQxAxC/DA8BsWiVbW2Hxb2RQ1TFcIQ0VBk3PKsYhM5sAZ88gj
7tbX2YUcba9ruVi//luRcz6x9BgJLNEntagnO5Rh09ciMD/s5HwE8ANya370qM6t3qxIN2b0W75U
po5726xkHJEg704KmoMyt7KZHFQCuoV9DelD10qeoy5bRcWaaowZ96TdqhBeXutao/3+ZVp7t/rv
/1YB7FqFmeR3/TwsmGna08YvU4WE6mUEOEg6zmqRBR+b3UHxrlmyfTRgjuxivhXHkAg68yvM6P/s
lVxI2x3dQJRI22Ee9tRyY9MW30iyk2SqrMhceq96Z2HIAwb+or4DjWEbBxqhD9byx4JWo5U9TFGz
iRo2IC2Xr9ngj9ZTqLxQGaemVx6Mx54xt7wrLmo0VZVjGC0miMLAAHKva/SeQU1ONPl5B+xnFP67
zHtYUtralbd8nmqpo3wU2aGr2MZKn/rrSkRLY4DubQLR1sifVycpg9Tnb44gXxwamE3riy2A2NjW
uVMgBiJLjhHGdlQGTivS5AKYSOt1107MPCTo1IaGvfE/rutgLAo9d9NybgMR4sOV0aoGUvBhCG+5
BDeowq5x7gnMhX+mEvYIT1KSbBU1AL9t9XilccLvstGxxmsKQpcS1unPJKBXcwKRJVakvlWbzQBI
obC5/WUnlV26IaOE+bu77m/Lj8qNfqhZyg3vxsytMgAfGJinCc40+vArmZwi3C5vy6wNcJzJ874h
eK2+mTGmEStVfvnxXF7o5+dzEH9tz5Wbt6s3hw2t5G/6+4l0AZEk4sy4VuVREpJ+6DZvfp8OzaHR
zQSqMItOxnGyVuDIczc0OyKP1axTnIGjOpvyFIVRkJX+ME+7ZX1rz+TOCb4HoVutal13l9AIpi1t
Bhig7tRJ7BcR68QOgML0pb6FxIP2wlZR14igFGxQW1YUQeUBkcgE+Ber9VYWzWinTgIXLOGnzrIp
DFe7haPAv/eWpgJ/A4nwt4JuhVo41COzf8gcCYcJsXnhedI5AL6rCHoZrIlps9d6JoJ6pL3fDkpj
VL4W56V/8t9z3e0EGhdQlksgQzgUSqW43v6ILwF30x500vLu88bw+Xy2ihKcrVbriaNIVOmYRpJ0
nn3/rH7XrxGv17U1o4UekVFAlq66a02F/9A5kBOEeOSmCGxGwRHYDFkBk2glH7eKs30jw0w9GYe4
qgYkc8pe7OOHSCGcLvFPeuSyyas5Sr6MJBR/Bjx0P6fgeWRSvegC4NDnKuXKnwozjYvynGp3pi7F
VvlXIBBWpNdekJY6LGAL2pRrZKl0OujdeX37nWqyrvK62CRUmq3keY4D0g2PtOv1fNuDe5ak2FVe
E+yMB5Xizz5a9id0S5hAT2dM1l0rc3rRNufYGrtL0WAs5eZSdPClh2OPwcs5dhaLEZlN4ueaVUG8
MPcyt0KfK7rnkWMnnWhlUBPEtq11yqapin3bbFjmkoZqpoN8QclwRrb7gzHBMnQAcim1Yuday4tv
RxXt8QzgKFlmwscnYJMMqK38EECerPpc7CkEY/FHJpBtKllmrLkRX3fFH9tBhpCPHRvr3bnYap+I
o19kf1TKHygBSk5rtkXQGL0E2NY2XvfFTujKcv71mdiFv1vXGGv8DW16+6s/HWa0UuHSeUmiLmx+
4W7YTttm9+IlQ9DcbGNTRdg7IEyZoI6WRr+CCvX4A41iKQNW8ukwdw/Vwe9oeaL7GZIUHXpvO8mS
f1Ao7EF6GKhQ7BWspel5An/40bznptz/rbOTYGPgmEugXQ3Sz1umv2Vw0TY3T7KN/4SfpOMViMlM
t9rztez7yLZZTV/eqgcq+vQGR8jur+fmq6K0Qjijd7MhnYqzbq84Wk03gcg95gfIrOQyjztPEfAt
3y5dgtwCwQirspTf2r/TuUaffbHxOCGDYfRzDJ5X/rHjq/eIlXVVrfryJY1+LPLDUtmfnxXN4B3n
BtDGxQYesz7CBcrPdkqnVYnU0aszIKoMR8ZWzmsu05I7ETMzhzniMeO5n7fJ1G9uzQOh72QJQqU3
T6oU+uTOjHsrurFAR+QpiQ/te6bYty/PToETZfKBo+VjK16DTFeRFY43kv5LEgRCyh6IBk+fkdcc
cAwpxjjZRgMvQ5AZ9hhFkaqakDrxyIC8T7lm9FuU1qA5WDtKCHx1YU7uWlntPLICoLJo0aarlM43
bgjFqb4X/dibTy5asogx4XYJOmm/DA57N8VJQAvNWkiTjUGrAykXE6Q0otlEpFYkT0duw+WNouCb
PQ9gW310I9wSm+HMzl2ZPf99VjFopWpXB+9uN72E5w6+Io7KDgSlIyJIsFKT9RCYxzMI9s7ogowl
oNsgIEHYrMB+1TDt/R8HpxN2JQcTjbIdoX3IJu7BR7UE4ybvP5HxdiY9fjoNErwP6RHJ0p8cMHIc
Hy6l+0u9eeaRRvCe8bZ8hJnwrB4yyvK1exFSbkNP7A5oMG4TVF10B1IChrvQNp4Uqch+nVwiKLt+
ZMVJ++9PC4jymQW0NsjN7AP64Z7JRrk9Ae0LLdu5rDDarOKH7UstCwfa463I+G/i4Lhgxaq1pmKl
ps2gv9WMZl/wGCn0qn/VLIK+asei2Ybs2LkVLp1Fv4SZqO4Bmh+YqEBvQvedEukAr6A13Szi5XEj
+8qOFvMGdjN/x9pnMFpR7fI56QLA9c32fWXnsPR50PbwIzE/i6o8nIVXh0l+JSxywIq/aiGsDt5y
EAGqn/80FaZAgkh6qL//MvGR0Erjrk5lOXp5pyVjmua+Z9y8RIRfHWpn1Bi3WZaGgK9u7t5RxblP
QMy+CFsmkNqXoBN4cbOXAC0fnvKiWkaTzVaYM6TMPAxjsr2uTXD6OApF9ktzAp7jza8kjcU3uPLD
lHpIP/py4ZrmAOwcTIfcF1XGje6wZyarTs6uziOpaXrfxt6hAYsOxWhIRhLlf8HhWjFnFI4J6H6V
WtE1E7xuiyrv1oDXoZGN/w+T9aJrNCI9+YPQJn+bN4Eez3LlntUT68peYz2P5G2obYOk2rrbYm/K
8cJKOUmgVdjhpGRwHem+JTi1Fo+ljnngrmT01PMiIDOAishKCMXZMcWlWaqjLCrOElXFIP2llFIx
3msBeov87X2XevIc+Vg7p4AdLcw5VGl2G3WnqXkmnYO7iWMs7dE1zBh2uXNT9kRYR+jOVjMhtjhO
tlPN418dCo6FgNNbUg0RRen7uv554oLlDo711A9XGQF9WjupE8Cd9K2RDO2+Y1SVSC2KQEChzLkA
zYTdoKsLgnt0wGxoBp2iB+vGub5aD5YvKtH5jsDtkeBjBH0VLYORDJRd8bO63qvenHrB3s6NIJgx
45t+SmWM5ylBKb/bN7k5RJAFDaojMJftBeFbEfwqry8osAaNSSNqJyXUe6v+2whVK77eQIUTWcYG
r+UCORun+9NzxrxOI+4QxLWHpHnqxHMnQ5d5CH7SaRmEgCPj7SpCwaE2WP/rEjJCjsawLuen0Suq
AZOE3GaUQXcj/zjIfchn3ia4XKnkKTKlwN9Air7cYBT4apJw4biEFlRnoU/0gaB0YHkOn0Pxr2ul
F0iOQOznzvCe2v95290JjdbS2M+pXVNZsnxbGwJ/bK+L3Uyh++0LqO8ASl+lfqK8v6jF6p3lKhql
dBLPjFaMU/i7BqxzHdp90uR7JPUQPck5/zomgoocfRrQ/2tWTY8Uqa3qKz2Qqd5u+SaiJSFeqxTl
6BhfJrGik0TTASKXAN3PRU1tvyEjUaPUgdALE41lED41S+xs/eBOkEYry7ZBmKj5paIIfcQGkmx8
6aENrIGFZuHjp8JjnbZzqsfiv2ST+pPIJQx6bPQCZXkYr/M86m/TVr5qRlveuKhrTytHm2UoyKLL
POWlLNqTrehUkXeUbdDrYfkj2lRDWURfxKjFUlDxVgbo0r385yoeOqoDJqobN+5jZU4w7/BNPmLg
hLCOubWHy/yf4HaRn4VFbeW6r0Lf+xdxRJ+SF/tMKL0SN5lOGKRL3kZapEswn3ib3RsKUzBsqOQx
tbjrI8LmHswubs6Xdwcm/giE9aKjNdxddsq1LIza4mT7Pfetv05HXMq1yn0F3PzJvGRnBgnGyLZz
8xAUrbzM5lwvK371684ctszdTh4NIiZcGG/L3A8ICTz2Q+KvPNU8+PU9zjFcDuVtR3npBKSjitSG
DbZEr9X4q8AFvJq7zbDt24WDIoMypFnOJlqy8iiTHgx51PCNr1LTZzFULZXbwDtDcv8HY3ptG6Vd
7jpPJX3tiif2gdgvET24G8m0kfN1TVYwHTYrG2blAY9QVbRHUlggsSSIwFVaN0IFqk1Dve0uBx9B
COnMJbbP/9GrMhXbmYhm7x5vfo3RSlWxX7eWdmU79XknPgHmGTDrBqYIASPCzwLHYl5h0SbzlQaH
mWM/wshTg2QSgbjf4O6GJRyq42aN5zgqRVwwKi9ylNquoxoQC3OmxF+dX79dAWkVGyw9mhkkuJur
2NJosZRnJLdkch8dvIkK79ohPNqii14QsRH0GiSLVg0A8+R74/kA5bbUm5bVKiO8pAnTC6CTGKIe
CoyUCCPoEFSPEFGoe7b5UoCZ2QdPW7nlOLocYuT/mNclZaL/6CKxCI8TNh0fLZXtaGtuULqirB1y
n/Qny94vjU+5TWVljrSdiQBlmjFON4qF5NGcwSjuDJJoSZeDzT+/Y/2K+y739Tr4UQnUEN+8tkyq
CANir380Bkinkj/aKMhi68rR58qM+s1fRZP9tUBTwr0Qtr+6EpTcUnigEJ5oVvnZCHHsM9zJ8O0v
N7l5K53/fz72j9iVvPJTKjJ9xdHpDypd6ImWf/RCITIgWvvJ0r77DJj4s3WZ7uIRO1jBayq39LYL
ElMuLdQpeOxXTM7pnndfyj4PLYANz7HK/puwnOTE/8Iyfj3aeoLEroyaxFmFVcVhHpsDrq92TJvI
msRyOTIg3tJUXc92CBgeLhYSsyyciVFtgpTzsIJgNx/rJgS4x2zANuck3pEnsI69gnjcZMsTTkam
ASo8QKFTG+iIezMIn2H3DXE6nucuEdb+pkN1iGupvDGLGAjYCR4zA6xY6ftAh9QM6hzNVtdzo7sr
ju24CpeJ7U2zM9SoZxnayzmXRbPgdbA840whasLsO1ZIVNNw6b3v34UIeco6d+NnLkicPOAMGtC+
XqXAjrMBk3rN4kp1hFUqRggYBhcr3ClRPMnQ3sUpbvvj6GAJgb+zqiCEltBhbf6UsgwOS/YNNvUD
RI5KKNjZYIEuxLtQY0u0ZP2l0IvKvHcLlGNTBsHL8rb5s0UHQpFdPvxKlAd+6Aw/J4s/Yx/3GOpF
XpS04iZTGOnGqP2v+Sbn7lb7bPgf2FWaRyJKk4w7Ez2E+rgqRtvmEIQTb62G0lrExtg8WPkRPbLc
4Jwj3qdfg53umU0LslGvAzC8XLmA//w3P40G4+1GsXMBeD+5rwP0yuO7248fI0JyGAW00S7c3PWt
RUgs0xVHYZUYs+0HII751/07RWTLcDVgx2AFAoyG4imOt0GYNQikj/gcUJaJEp3uPe/SuJLRPhrA
u3V8FjS7eZZ9lB4rdhtvBwkpR3/dZ2ncuMLiycjJM7p4GW2iLnjzwRoLBAR/wl58/cR0ZnNeCE0P
emin4fY6eMXhO/IWYVPSdFDgFbEBSvn0NuMRqrxcfwTmYlVjbCmoibha1SVLnrHMi+QCH1Wwh9mi
TrZJJSTcvFssBqd5ljlP+EYC05HXVk2IocHnrlYtKSAhgxomE/WINAZYXlztkow4R/Fzt+9vZQDk
0BNYNPMgIlsLNEAsKERzhd9TC0UxHLxrcB4uPgGY6hWw+3KQUR5aNd/cgcDQHuY3l0bHcUUDx5V4
s+i3QkRksV1CqL79uspp43FwiwZPRcocE9jwCNrYyJDzxvXWch1/ExSlSBslgzJRUx/i1YAGFSlj
BEXT7ySmxAITB39MtU57emK0sKjcAPPApHk4o2704V+/psp1cF5/vNof3adD/YQ7A3uf9JBSWWMp
sIlXupJ1W3cVydIF3MQHNV2UOygXFC/2YhL469nqvjsksOJjy+3vvnAuFnhvUz58INyuqYUFn6HL
EBzSvZCelUThK6PBZoACifzKo/nJMHW1vXzTJj9PbK8wbBXronVXBHYTVXmPKMqUxMo+ZoBil/AK
nMhwq00cqJWqYwxKqrSkimrp8p4Erme5wVBCKyHTH/5HSwSPGAMGCAkww2+pcw3X/70VixPPv9Jg
UFp6SDeI5CS/BsE+h1XRwakKaOt2sgjaTicLfJuwkDx5HEvYZA4+5AeG0OItil3GDZWhXVnUWCie
msRWtHN7+8K9hlVBPKdDDAvROKXYr83hZLTTl/bztEDT7NU8pTafSfBQc9i/vxMQEXpRTwbQG+K5
YRHO32mFtEJS6cZfY96a8v+xbd5N4qTygI32IKDZIq6d+fyeVc0Q6g/5633c+nco1xtX38ZuUCxQ
mG2lJ0air91qcEAPboPm6ge6J4UHlpTq3VerMYPR4HSl++yG6kX97eg2sfF1UlXM5FjUBjkYBu9f
EbyOUW2WMIrHOuuInpbR706DPRSCA9Yrt4XNTCAcLDtY7QcxlI6gmqN9IMgenjmRABB0mMoLwdar
okl20/vDEj5sJz3UeUbDKFOT62llQ7mHw+dVzk+e9bqEgdB99TEoquotYSWzklcSaDjsFs9KD31q
nZnTSB67MmJWdpEWAM6am2j5cyrDR1ERqW4MUZghaFmj9TRG1e5GmK4vfgekCv720UWTcz1Ep4Ra
RkbJKVNRkqA2ex+AGKP1j/n+2mYeQ1jd1lWcA8hN35UgLS32UwBBj2bdrouFTDACerBUsyDLHvsy
MjrtdcQWtvyVD5IvZk2WV+Eq+B/p8Dsv3FeTO52fQCxI8EuGrzNVCKyd/G7gYgFmc61FRtmUVceQ
VhagJrFpR3wvAaS1y9Ov5e9VE5jTF1Tbtm50LECheTw3dyMjXw0J3Mrv6QxWYdXhwrzKKrt2oTEv
M17GMKeg7JQ55jvT03vnAS9Hhp2HkMb/wRk742cNJTyQWcVesErRnmSZ2nosm3oBJ3df36FiotUg
M1Y2jhKqJlz01OK6sF4YowLVCq+KaRRekbBZIZDGu+0szx/pjjYugUJrCz602jdfJ0lNGkmhHzyD
Wz7e9GA233drzOv3AF0TkTrTXGkSjhY28+JzlOc8VJmD9GoWZEe877ZtQHjldJHXebMLlWXsgFl1
4Amox72muDo/VHjG/jpc7k10TGHtE/LJoLA24ZGoBPbZnkC/W15cc6oYXQFFvIvi5X236PI7MQ8Z
99I9598HyOIl3RkyIHgllEc0ATld6khXDOBGHJb9k1/hmcUG7q2BiA4bxIver5o4VaC4q+lhNLCg
s9lbKL3G6hMetfjPWpqbGaHPgsJsci4TWBIqi+7GbCOJJsxxwdkXPrp9gJb6yBbh8Le9P5FGio9W
xS9wuVtfNZvJCC67xzqUII0ObXOyl74D5BhidtLXF+1ypXRviEcwZcAARAGA2ndHcBdySrR7uwbf
mNUYKxUQukmQDAa3BXL/B+VYSJGgntsL3FeaZHXOx12d3zml9Okqbbm3x2N+VzgxAqBplPhfMYAM
XlewD3KiZn2Ha95C+YRI+O9VFDYh0walDm0DrMU+AWmjipfA8eLMtXFxBpokUWilB+kQrwsqgJZ2
LUKwMYt+hySHKReLcLdcDBDT2Fm8wRpgfG1zOo97FTsH7RvxBp7xFzL1XtN4AwhzXS47oWaiGphD
S37nbz/9jZjUFtuYe3gkq+q2dFXAMjQ2tnNjTHrPlu4WOdkeOfFQ/3HcLSaYcA7hBc8Up+x5oWCR
OgQIINZl+Os7v+7Dlr8pBWmFnZFobq3yQ9bNdrQP+9MXEinxorlW9FI7wJy9I/7f/61wXFN6BUz5
2GqO5idMjB6iOC88H9e1KSS6IpaicIaVeZk2ibnFInwOerARumhVrbjrN6zmlDLNBvDrKMY5Gvqj
KkIM6MFM5DYVWkoVbTo2Tf40ezWDFoFPEfAcyFaYi7ctRZ48p97l08NWwTLfv8eoVxSgMiFbXoFs
plsrlV8R35nKoPuXip8ZdsIdCVTXoIPjK4NvoZqYCu5f3nGlsE46J55sEzFNKrH6Iw+MMwZclob6
d9rcqLSpiHwLGMsPCruwn7m7CsDfgJLQQS0Fnj32ZBJNZ+DPHwZL5149GIdj7Oz9RbKAf4VVR4gZ
mCVj+V9vCQeWghXMY7aMPvzU3vPY1tzmxFTLCR14YNjUfSEzBjAi6KXhIZ8wHfxln1Rc2PcUdWFZ
MrPUd7Khg2qa4VfAqZ6gXy/EzMtdoBB5kv3WaD876Q0cn4Ixva6D+RZvBC/Zx/6OJddGqtUQzYat
DQ9l+Zb+4Jdvr5q2H0kRys9WQwOvRurcthNwxTLqo1BzLCffZSn9ryOgwg73PPEgp3ANykEtV2j5
ktdU8WXVHD7WKi2H7QrwMjxcXtjAW+qCi8JhUWOofRcdt8V5vq8WE1SGhgE31Aqo84k9w+xbAXe6
Cl/SnRmHwPaRf0CFsitUr8rUxWCpsvewuWJpe0Q3UvLkkXAezLG0b5IcClzL3eWEkKCv3NN6t3vB
bkcRDDCSkOtTxUMsp6wXKoSed8AbVGBiZqHnQWyHwmMF+E1bFmm8IuGto2Al51BAbQIGgYXShfQd
ut/C2zk+qNlQiAWHBbOLL3BAeRhGLUX9Mr6ttcscbS0xZHtpFRfT6Sb6KewogZ03OliToYFwUNXN
sthtDrQh/OLpL/juXsZfEUt3rqAsZptHFKAIusvhXK9+ye00s8AHhWaER/1Bgo2Mjg8Yl4YrQoQl
WAMHSMqtdmYWKNN4RvgcCGcBURKvV6O/01HsnwA21UI/iJ38a7ma411wYa6AUpHA0ebof4L2g/VK
znaEED8DsBUcfEKmIxyaSt8prsqZRTYgzU5Ut18AaeUyEZzTmQtuHE65lxeHJhewhcVSPFM13V3s
FRoBFCB/rYnswlfgQF8oNIaW0rx+AJzY271jKUyYxTbeFZLPp6JAhDJQd1bM2eqOwem+rcU4PV82
I5/kAsAAc9bidmJbWCqhg71IIhG/RAcKMnhHD0KF9HWvk/NeY2TwWaBz1S2qMmdw1IC2N08TSEQ5
XnnqBt51OQoU+cQnTx+HSdw/dK5+2geLpiEMKETsTH1J1ajH79DXTHClIq0IVownUZyP5uV7ZQbl
Ix9f74vfnvJ0RPUJgK6m1BGmwWWhiXqgxDM6TrViBpQp9lYgjohBBLzylJFEoCNgGTSlL4FWrcxS
D9VhF20Hi5P4dYHs3tNci4/1al9+IRkWnngbSe63qCd9KkOzm7Xt1RhmsggvHTLBS86zvdZmSnEG
5t2fK1RWMENGO9YmTDjC6IvcZtFEFrpSGET4demFyPuV77Am7dgoJ/1wqwqw/inpeS1A/1ie1+/c
Z0nJHdjbeUzfIPqO1lnpdh/vEKX72U3mO4xrdc1MDNrBBYrMn7G2bnA3bUiRXCSVf2X+PvXc87Et
wdBtWXyYRxjDA1xNVtESuY2/SR2tCc9BYEKy8fUuPB1jdEWSmHfMtSESZQMvQ1XhdVQH8p4i21+r
1xoKaTGishkIHN2+kIHIAip3sCohFdj6MzNxC0LJbnjRlZPF6ceUaSyOOCepjs4giTRsNXNmG8Lm
qKnVqmSEGqpwvYAVTJBYya/vLYkH5FhoKNL4rBAjuMZT8AEGzDq3L8XQ6gnlNm2dA0kkd3QoVlos
FGB2ZZBB6jq1rLQLV7TUt7PYHohgOGwdkHDTrlNW7K4ympMSgxgQyD52ZGzuBOggr/wgGhopZQwq
YeEcU/fc4HqqrIQe3/wRtv7bcDNMAQmnk1NIqq9ysG/LUbokg7JVYpwKdSo+9xs7Ei6VaSj38MrE
GwPZYzURREDciJk0RA5Te3P3YuuTGAoJzUpY3hmM8gFLDPOxXz/Rkbd4ZKJwzfmkUMcWxYlnNh06
ojEMVUiVGmJ3S0L3vpuVLn9r9jz+eUfdqSMabjBZ3rd+3XFNvL5TMswTW9TCgYsTI/zRqExn3I5I
hNzZJ5dP+y5d1VoySUhTmiO/0vtvzX4+jum9Xar9iiyw97uLFeXmF4Wmm9LAppZ3c6771tLtT7B5
FcaopYZZNlSkanz1Gy9CLtGnOiXW6tNG4aCyKGJ261/KfUWKkdFc3g4kSO2CuyZqh0T2jf8wOUgN
efHPsVrvS7PBcGqOoT6UjlK7C05/v3JuB1KczuL70mNkjgpnkfUhPQWKeajQ7PTnMbeLgp24DDba
B+GtxImLvSBLo89CQ29imdA6lC4W7y7YbL02eNYu/25qiZfVLipJ9YxXEXZbbcWo85PRd2Yid7mN
WjbwbHu53RtxrFFaFXmKEyGAiqOIv65ZU7oEzgruCtnqQMBHK1UjhSTiNanpKN6yvEy4gN5ODIng
7hHF4CwQnjClV/b7IQJmIm5PXmYk86NswPSCDuPihiOt60UasMTIz83p2+lSXkWf2UntKtCsBjdY
f0qgvFPlYf2BE7sVun9eRePTln2TVK/tMrUm8gjMB19YtQxGFX1w+yb6Z//sk368B1WEuGUQ0l/3
jOGq8z01RhURQ2jMd4763pl4VeAhvdq0THVH1qbax7K7wgcPUTZvsA0fnce9tKrlTzNmE79h7pw4
IR6Jd3fa0L6vk+DeFDnOufY8oLTqj3+2h9ZGC0GtAPn9QrlZxhCrlQ2s1fePz8uJG53YAsg2hGou
XxbhH5njc3mG2v5swMKlPLKCPsTYdyaL84pUN0Z9j7PEqhUd0QErGDgg+EPml1D023ndyRp/khW7
uAbTo0YG6mFtvsbn/i9w8kQAsRo8Y0ZjRNj7iEP+vFzs2714Dku372I3I6IBSGSU+Dd5CQ1iQYzp
aTvtEYXZH126SBdBRvvfFEHWF1PTF8Km66zJqi090UGVAiC+Ax//aTZrEBs4SmaOUg/hVkfPySbA
VLdkzW2+4bG2ve91mpnh5Oyozw91uWIiK3oX0oA0g1sEKZZra3eWVzydl0HHmZhYkiEENNf2oDdY
obgVVgYfAQ4fz4gfCyFeloqkpOCEjFoHRKQsnUwiD+h24SYuQ1/C5ucCxBxCrcXQ8XmLJsssBBcR
J12ybkZdwutyaOPuPeX8jRLLh0nJNzv3CLef4K6KW/F7dG8ZA/obAa5eX12k2ui9Q2tIRgGbvhRh
t1Icn8UkRsckPS+KNWlEO9JhxqrPNUPMRPJFGnpTkix2KUHJJm/TO/kDZ8pufqIRCXC9UhGJ6YgG
aKhKoH8eGkUs16NtHRrgby/9DQ/NVjxEfbxKrwN3aAGTG1uQD3ZyG/4GciNQSQjedqosaRWbi2hy
q9r1XCttCgv04HGMKB9Aa42lKCTcYffO35KVqWVFjEPmJgwZ1yPfAvKMfKqwC4T0pwatfTBKD1aR
0+PDjvfiisxV4lXK3MpdYRnsNEJJYRNIDqeQ5tRtvZ2wWe6LdIt7J/H5OHaO3jLIlJ9T5zJF5Gys
QTl5jfW6A0P/1SY9LrvdTCZlxRjqEHBIAO9mvQFcMsukTkunR8mkyXTKbLBUY8rK5+LWnzRLCME+
sog2qhGGGWmcGecvB4td0k0R/gHXRr4P3Fu3vGxP9jkagxk5+d4nVV18fPWwwIpiG+zsoOP+c2kh
HJWhpXM6QfdKEcikAoAi/Hc1rgbDpcfn0ySJhpEiXq1jVTmcL5Z2L/bF2IkGnH12JSW+SU6Z7wLG
x2HXpp5FuGVA3C8nsCz920/vw372JccSDIS7n6pnqCC8Am/613z/dtpLhr7t/1NkNec+KhRpDq4v
KVpsa6EgdkygKtBwwJM7imAbdC2QW7YwlAdx3y7SiT1TsYBJAvnd1grHg4e2kN9qtdWkmOMtxB81
2ce3LUbOijhgggGJ4V5RbV0Bm+yRvw1IkZTWBnPHN3Cr4RJTGYCMa0dyFAMhj4J20Iz4OF5c1Wk2
yNhxpi4LMuxA2lf4B11z0PHtCJWJ8CcnVGP/dLDJygkpIpczdICnZkzkYl1ASV00HvG0Mve837OI
BJEp4cDgkEBeLLoFix1HmHNggZPELiQg5A1f3Y01DyEVNpDWcf+oDm5NefxL/ywN8M4DuT1K5bzm
xPw+YiTmFkg1M3WTE0uh9Oi2J6IMGO6O7Y6+LlP/Lz4xQDCDHOnGfiuNBX1IfW9wXqLyM2H0guSP
sooCIi1J2YE5TY9FLF517b4PpsY/N5nwUznzuA3jcjFyesDOT4VNRSeFndj/e52RP8cxH6pS6dC6
PXHsKsavXjGquXqKipIYUKjfQxFQlkUas1kUrj/9e+pZSMpCfHJi+o+H3aLB+tvxO8GM7WT6H56u
B1ZX67qreICpnQPKGPO2k6Tql9V2Mb8r982dSpY2C1ThiM/rI/pPcWMILlJF1TL/Ad0/EAltDySa
mW+GjtqGksrDbLOoQxQEEjPkzAQLgRA3pj+ha6OEqJOcR9iHziV7oZZZ9wOriUyTncLubUf3h9tn
41yRCijidCG4xULNpg4l5eIpfAK4jAqyTWgMt9C1bLgki7HJh6JuznOFqICBcvU1dLptIvurY3ot
RGHFvCmfzyloGZwG60BbFf/cPT+Kr170z4yvDDvuuMHDc9RHz8sd8J9gRXDHnE8T+FhTbb2nn42q
kBJEnV4QsRAJBKpS66dWHBb+0Dtll2Z+SPHInniyiDcFXZtQIehcuWALVXgUUAVsfyCIHfdlPWoN
3fAJPXvnndt3qHQ7fGWXA2mGnkpOnt/bwy1EHCRqfiaOxLFa44du7amrHBY05jaxXPS6Dll7ZALn
T9URCzGRyRQ6tWq4xUokH8H4nXdDAlKxUCc0disei0csmG0efGrNdQtvGsXz3oQ8AfVUHPDL2q6O
jXq03Q33jUNuTcuYysilRQg3mJsfMoinyJcyrf7RxEMU6MeCYAZom8Hvyvg3VubrIxBbItAeBLCK
vYMIW80q9Vde0XPs2Jy6B9XK1Y/YdamBPvmHIX5Fjw8DyMrAYouFfP+vi4z850feyksFVfX/LuL1
hhFsMzoWifmKFwfgsWLCaEHYjaOEAmqqLF18Zj8zBkybgLMvntod9QJJ1DZp7XKLxjKu2TnrZJZs
XtTzU0RFAOM7z+I3KwYeDb0EYWnIpckySMsFPqt7bRK1/nccY9SeiayVYrl+VEuyMXIEfjX6fHXQ
+ndjTi2BKIxQrLQYQ/u3QbeG+GN5bCkxAadJzFX44Mzl7pTUQMOv0+2NZqh5j2KnUBw/WI+ypOcL
y9ibmtRja/JA51pHqI+STBOJP0gelZmS7fM0IsQtQJqdfyCaVnl+3l408HhOOUphmss534RgT4yz
6pRv0wp/oNmn5ONZTfl8SzAmRiPaJQXYExsX/aK1WYKqXpz5TkXB5xn3ixzHRJE5pG0ue/cBPfzx
pZLXKQjFq5yZNRlf6f6tgTKb3NfO+hzeZFqEOiBSacYLA5BLTqYH1i9EWoEQ+MgZRiY7LdxOph7T
8H/5CW3h32yayga1QFv5qkeumnnUhc1svkOWV5UQtYp5Mb+zcNTb9LMuVjxmLnJPrM7oFn0Gqu93
+uCsmLztvyGhrb3nt7AnBHsw6iseaaqkMx4WBql3Oz19bMM7ykgk1j9s1jTqzQ+Xa7RVf64Sesea
2WVY956ukHH5RYQnj7iDZdJ3962Brt7Hj8pUYzm1aULqG+Ma7d19aJdfYMgnGQE1gaZ4qJpBU612
YQ45O578mdHWzsE0k+Qj37Hdzyy+/E5z9hLH2sAFGHcS9YztZ424fk3hmEKgVX6Io96q8gyGvckR
CC9XnrLknnU8krWJYjaQzybRliSjAJbTuLjdpRrdlfxRIz8rr6suT6T5Ht3jlCnEHEg9mKqOzBp3
SwlKBSfuOFYj0pEYVJKykaoQiGM6ohWwzWcghqFE0RnOrOstMluPIf2WYbxBsSlKmy47rmFlueFn
9YgNXwHPBnBaRLhcWzQu1KSy2bK0IRIivUsl6Z0ILwDMvqI+gCvJMKuOfPfJb7rswZ0O4axExjgn
imnXP7qp/91zj4IgBrj6VBALmzgcOnMZzHFT6wQ5A3bP0jLOYor+pbA4pJ6Sj2/yxGXnLZCiDngT
ZabcGxKRuTS6NVLfq/l6fEvTDt3nUh3pmubceHUmvdahSJJ76TepyDcMnuKlRV+x6tnx2HAqeN38
vmq59hKqqsHpq24w0BEyei4VE0HFMLX0Rr0hhLPDBbzhQ2yDpM5AzcZUi30eW3w2eUK08jTWoNW7
8KGMo18zpmO4+N4xWzX14ZKn+Q6yVs04+dFN7rc6QoLe9+2ooIM/x8rb0ewwJrl1gCNc4ZWb+e5J
qu54UoRelxd2WZvmI8OdNBxQUwT4ckSTH/2Mz8iEcl90dHrv0qYGOv9A8XMW217cB8ZrS1e2wDwi
i57siFjeEWVaatLejxY4r8D53WTh7ttYccYkUI/DugQJYBtH5WlhLOfvvMEz44UibzJ9y17K1YF3
wMtI3pCFVK2zmrDexr2+BEuAE2ADdbVUEYXhGoJ1CKmbNmTXa1Rd6fhs2KMcXoPbxyFUzXvr/ABk
6oppaxldAjT4/YqGzoq/JLgO6UTsdpAjlLiHFj3PuLIYPZUK9pPEXnPZ4AbKgIcd7Di2zzRBI38A
dXrGUb4VetaPDxGWX2GrLvvvoN3LmW0TMJAHi7ntGSs1CCGDaovLVbebMwHX+r/VpnsS5fYMyCZb
SLQFPh93pCdxFEMKnJFfHocYU04CgcRy1eaIvNXZsJIWvDqtrmLl4zXFWo/BVN/3IClCWTgxe5T4
gxo2+TBiWPhWZoBFYt06Sq33d7GZtQDgJTY0gPJnWw1vHbczGww11le5qPPE7VBRTT+ii/GOMpMH
O0wmsXD/fjkt5ABH6wLNCEkT6oldpwS7wzcTjQpieuyy6n05pVDIrJv623ZAbnKXCFvlDlwiEJXD
VTyL4CgMn/SCovxn3fE1p0TjtMgjGPzUQtmsipUoXZg6sE4t9UkPQzk9uW50/EbZg0Kdb56SRXU3
32XhnZb16bZvDl5PBDawYMxNLnB+JYvJBJaL84CdPvKJ37RM+qo92ZsEGQVIVR4VsNKoYcp+FjBV
3IUB8zhCYEFoi1t3ukK6AwLHos5lVIk/QAIwd24cFTglwkiUM7Diyp2+MBq/3cJq/tAAczNZ7UmQ
27Phoduor5+tMfjlQO1cJez4Ln0ZJIcRVGiEzf+uh01WqZ9a5LxRX5GUi1tx1WaeQpFc3a++1v9z
wM0B6DCh2ge+Z6IEViaXfOwehfGPBvlEdE+OF4kE5SIPyN+ipxZsD27XP+PnzvDHs7m/nkmv1+kE
vdQxCmsrgS2FAjuYSK5AgAs+QLbARHGi/J6WxgiTym8tmakvSkozysk/yyNgLDS0lxNzCarsmrmF
fnDsYP96+6irlcbTERbpi7wYucvL4LAQBR1aT0qx8rC/Uhm54nYcndtQMlVrUIenn7eZugLY37BO
R5xLWHr0qY/NGElmtDN/O/qan3eai5IebbhzPMdln5aOlXBPiEOnpeuHqnS+DyWxW/y64AuGPHjs
9+BHuc02I9lsUC3Gpzr56QMgU1s7IptBnv3VXrGzIdtT8+DM+ftroA04QrMcc/3qlLL3j/oRzGS1
Br092dt8hvE4DbJMyutttmGD1mouyUPIASvIqwqwwDkQP069NkMLavQOI40WYHa3RXy2+onsXnIP
3DhVWYSHkdb1FuCmihu5yDocAFYDTNp59jxgDr1Jv9ZgHC73GPybL5nRyqlPIEyKOmPQ+D5mP6KN
IQDRjLNyqJIZwdOYSd34tcf57Es5K2rGGGNLiQkPmK4MmzUoxu7H9iVL9djD4EN8wd40u/2R1ZB8
i7+pmCZBZBL9hMUxf3KnOtj+1SNNEC+rTIduATFBhLjEOEyP5XGkJGQBNASvr2BJoiOXUHy7LJEf
PbztIZ8oy3BjKadznEdLKLIbrLfWneCIcOOgj5O76e8//dFEiYC3dhUGmSoH/VDrCREWFoDxW7qv
Wt2XVwbViZ3yMOBOeVBltWVgC9ttMt0x30n2VNiEFXs88uZkoWqg4vEnUMZ42M+7ng4TRwNfNrl8
L3toj1okL67satb8sNXCNXbqAymjAEwEWncyOiBDlDuWG1YBfBwxzYyOxejaOMkb/mI99J7RkHQd
CpwcuGm1DJ8dvAOOlvQGDIjbIFQChDfMoablYCI8umq0HXKxVptn8aYqNP3z5n0b+BWLVibCGFC2
CENvK9n3QGpvejPXKnNuCi0LYIaoojODZycJ6wOmhSNN+81yeVBP0BA1+sRqBr90YkcAhkcRiASe
rJaYMdhHVddFAIKJkEMhiRsW25z3oPrnv0Me2LHzGyDv3BDzKOmXjbqKafxp88Vphs5FbSA0ktR2
bOzz759Z3uPSdittx7M7vZ/nuczir4Sk1FpD63/XDlID9BR3qiThueQsJ3MthNGt4ajK4SF3EfXu
7VU2cjv5cLwQb4LKeo2NfCNvjPFQ5NHf9b1mIE7z3Sl4dOmLgjdGxgffE46Z5NHr395F+fES8daW
ew4p2Pr/HgiJA+WcDk+KdxxlMZgWJ8XSfOwfGhXBK4wyIMMnZRncwIBlK6lZIgAIdE8YJzHClpsr
U+HIZbmZ82p1bD795BgvMGMjvcGBct7Y1PdxeGz45uNVMpo0gXauMV4s2cUZYsRJYcFMrNxr+WhW
l6JdylVys9HWRYrgkLF+SxrQ1DKaAHWGO3z64oRfA4n2OEz1Fgv7I/j/gjok6s0m7a9kth4al0eX
GB7nYlZyvODN7JvEI4Fvlm/umVJfOZc61wj/c6XwCeUM+4q/qkuX1M8bq24u1VCRUgxicmnE6iby
4Fv8xGr/+P1+y6Ju589g5mrPuq2xzpujD+Cw8vmqrIdcGY9Q6AYrv2hGYw1bsni+SulU3mEANEKv
Pi+jH4frO0o1/kaOoNKzJM415XTKqAerXR44l01bnSND1D2H3B3xqyCj8vtT5EHIhoYOKj1EzDQW
NW1FItyhZ+t4ujEkVNxEWy07lWStbD9+shi0yX8lKjTrFiMJQUuy0WQn4n9wAPLi1nHfWVJqPM3b
BCTzned8vlq2v0QJXKxVMvf4Zd1MrLZU6GWfG1SKtkmIz/0NHoornrYRJZslw+rIncutu5SSFtAj
NI44XF2HVt2w9jkk96FQOmwIKb0ZPTqMk6WA3J2MeO2ZOe6xsfUAZPirFRK/EAovpFdLO7ndk5eE
8n5jg8KoW/TFhe0GGnlXiY3UGhmBpRnRHN+Xk6lCw1hl+zBAEG91WmYFYjS7ZG9aIelccQp/SC2x
FShfo2wkjAhacUSgBl8jJTDUCJeyzC2KZMxbNTGbd9I+cVLfF6MykhjcJsEp0Npqvbo84NZCCLwp
mKOrJcMK6LKrK3QwnGWV+Yw3xfJWKQZMxIZhTg/RoqFpdZlkOyVvt+hh8fpaDlPtDOAB78VcZVaS
3LyCtQxjaqPuKZPY0iJUDq66vlWhph5PA/xsUC6216EgBTphWT3lOLw8RlIy/8E8g6zamlehNdEP
o41uk/KsgTudf+wr/sNvK6uagZ4md/2vtxRnrdjn08Tw4r1QVaS03k9KizrxyuRjgI7L1P08u+6Z
VJO4rbe3omHUooz0j/JJwB7gIHt8tSidgJ3/6NQmaMkb+vmtlAanlGImbPMfC3LlA8jtqlw/jep+
elWwzCeRuRiX91/uSHWdJsWL9XopdtM8gTeH6cd605XHHuVs3C1dzJHNKY9myC5E01UXVDrpxMQi
wyWMRotAHW4MVJTuoc9XrOlRO/VR3rbSDs1POY++pGCZvAoYRmlGrYHqzrF6a/dYtWJg+UYUemE7
9OgKFbTsDTNLrJ3pBsBtjtS5fFH4lLUw16vMd4dQ1HxN5Za5kAUyyq2L59qJtVUZwAKQ/shQ8dTc
ohPxyxkm5yRVLCqosfMl1PoRzbRSF5InEcDNY9dq+afL58+J74dp00/WMELJqG4uZuLDJNTMMdX2
K9O99WLgF7L1gPNcx0mdHEz9PvJor6thUvPn2oOdOc22NQG8F+lCKOfY6lf5leEBKIp8Zouok1nq
gjchKoJ5DSJz9hV/N1tKfBp0XtLuvq+X1xrbnLDEYmfadViL2DA0CZ61JxLsy/44RmsSPPwe3pXj
HzCM+oNhBLjfrf6WCdhZdKeNvxJkAgYFHWbS4yDcFJUN3XfMoiVn1MJOju/pE7UreTAq4KvRYa58
76ydrhJwbhWf1tCqRk2v6xSC1FTRoBNhsFttyk3LoedTyu6RtjkWh6FjEHtHhXLUKW9f5ddr5BtU
0S3ZIUGgoMmKA5GHRX9d1AXrx9xiSuYbVMByu00frrgiQ5Wgudju7lPF0s/b7IulN8J/ATUAAL1T
wnouwF/8nxKgm1eBNzYAHmUsSqT5FifAA+JYAeXCA/frmhI4lfuN8Ob5p42Cs73HDChRqO6SqAbS
JEkjFdaA2SuPxS1WtVJS3ZLBrh6yHKq2UO+DXogunxGTcaE4oHLy4if+woFgVoWU3Vn5LDuiWdfr
6sHuG+Jvhf6r4LPa3GyDScqvtD983PK4vuuuTNVhm9B5gUt8NWfQB8N5pt6P5bzcovh5iUSQnTs6
nfRoTY32xlW1nzG8z6G2Wn/Bq3liZwFjF6xuTJXkCTQ4XCfFltthElgN65bQg8oN1FOTKAIUorFO
a65JcvmBCcmG/cx6ZrgLBdhQ1oMF+Q1wkDnXy1TZZp6NygKVsc20GVRn2n7uvDPWL56Em2XcgRr+
xITNkqaQY+ue0ugn/iz8RDTcFFjb/v6ew8NGimE/QyHH/TZnkiYH8K3ntT8W+BblNRwyMoDLKcqC
/A9prFiRrspVQSsin6w/H213wXSUP93tw8eXqZIjGB+otjRrsYV6jPh0M8CiSA8CaeAjBX2hk/4M
pBBDW8YKeR5TExT/fJ9tLqC0lgAQm6zXT5689jkWzr8inJsNcEG3o4GHeMtKM7q6GvcxYfm7377o
SDcLwsZzEXK9J4kYRFj6UrX98BnM8Q6p/t5LBs5eX4gIgEmZ5hIcp6np/U7x9x6F99vJZQoAM50K
0S4Z+Yu8U+jVGh7GhdiDoxR2AMqGQjhEvxogCfaCeYQ1zcXI11jcpNEzEOhkj3qGPRDY6Lrph8je
IKTAvpi6Rk7Z798XbXG2YxcDOermGwviYH7N5FCp1Ibux2wkCwwS5kzxh/C/xTFVVFErBs1P3pIj
4DXRYYQnGojEdd4QrQz5hz5+8j7YkaD3lme5+SD2T8v1G8vAz0bRQHyMFKbeNB7LqWzgY3Un3hYR
RUgMOo/5GbnrHeIw/IYHgnxOhvFkeiW7kmLQ4AnxtLHfjQEOIQ5VpThk21D3A0nH/fXFSBRlmpjM
yhaQrQMKimmGWr5d1Uu/7hzfzfRHt+q0+q/nUfRCCSK+r/luBIvAvJ80ujpm3v/qxxSW5SllfZ4m
jtXRJiGqZQs0EF1O6pinxF3gcJIdNsJ1pOgnqZxRkVwdUHCMQx2y6ZOSPUioBZOwBzxVIoo2lZJE
sj1SR6KV3581tDz5UuMZU0+0mTaxzGo4DNQTbyFVSlLt2vAAEXhLWgUry0Zd6fuF8u5SgDyZ82hm
taRu0FuJ5ELblhWMrCMaTjFX1Sm1QVkNGX9z1VrnRdyCjVpUPl8pE203PHW0qHR0ALOfao9FSa3O
MZb9NsHE2XJi9RmSuP3JZq7j2IKm7FYupED5fJGqJglmhfZu758VRea/PpWQLmn7OKx1x+k3arBD
DQceI4TgkWO2+m/UnBRVYeCL4oPMlL34UltzWadxdxdPvXk3Jady09KNosFpesLhs1aHSszG2NKA
ydlO7MNXQSDssw5IWgycWlwt/s17G/QrkjKwp3cG/ufcPTK7p/Ym6im1q7t5pbctTO6mzXvhLA2y
OzHyckqzDXxIA85ZeJ+OjpULm7bK/nhL4tLm3yYRCTSIj44VM6PgwzLc1ZGeOOxL8/1p3EcxUyHi
OoowLsRjxW+Hc2yANG1a2F6T48ylYtTJk972IvFgaGP+x9k/PVB/T7jEhAX89ejp2965yXH+mNNO
61OAeNqUHDI33hV6P3+kP78y6YRuM0L5vWcvDi/wfaSlRqMC31bqiDH628CrhXusZO84NsfuPouE
UBy75rYSxQ7UujM/TrE9dlpJ6cJZccco0pf3t+W/9UAse00VdmLEFtedjP8SP8iPU/StkXAW7LF2
syoirx7KnPQ9LDaw24cFqSUpSCA0lvq+ElBpf8htIWWK42clD+aCRG9Lh26Ga1eV/8f3LAfrjDo4
7D0LEQYI3EG6Gzsa2UZNwxAO2uWXmpVSu9ZTjNKq5pz6UAX3AfElTl9yuY9MSjFn/nuDAicfv6kA
bi1OKK1yi6x8WKca04TXv9fasqnajllE1Ecy2g1q2NEsAHykOnC5irRYOHm95XvuI8gyH5Ojx0dv
wyJWsVR2AWNk15GMSoWoCoSsI38ZMu7Hz+3ZJ4QL1qBK026dLCKwIOmeev4vmTjWhim93h9OCFzN
XXKtzbeVtj37txtGpDw+bvdRqenQGTFon7Ah50cOmF3CHXIb8R6VSyhY7mkjCd7G8A+gfDphv1zo
N1ckpUhz67PQLNw9O6Eg6a0A5tMrdjBH1hDeIxATzfkhgSONRwwTkwntLU+UvWqBG476VbqN9Z2N
6lX4N2fXEM9/0SduAmagYbv4AW4un/sewvdanDF+g7Xoga6BNZPiX2emDH5zGjwpX0wNVWPQPGsQ
lhdny+23Qz8WYnewelgRHEC0zsgN2Va3SWQTJDtEpplY2uBpSclNTI3w9quIGD7zH795PwldMLel
F/DIs2A/T8wB3C9+syPY/ZqAvdVpi9MFJklSTpo1JballJp+GZunnOqWQ6nwU7BggVLl61ZfroY/
raI8xyWC0aX7NhvpeR+27nwElemN0hEyVnOUTGiosuMygpV6dBpbW0yar1pCjqsd8U+DsgsAlqto
BCxXVOVV0lvs/q35fHOT/Vz33VUNjz5qcFGUF5FeCDWLsXR7y82xrPJET5j8bwEQV65pjrPJ7qyw
iQ3OdEHw47ucOuq7M39wuXA1gq1SWfcxW3F9zLgox8ci5hJfVayYPh8QYA7XirIroCd/OaXTzwhm
W0xeL2U8OOToqCzKiC5voqHWMYpBZPGZPBHPBq1iCnS5mNK8Z/ISUc7XYoDUWYs0vCqh+R5XfTJ6
KnSUFLEF5OVrzP3tbT1+hrph41m0CRxnjWLN4n7Ih5KAyy+uWcyk3yEXIb/KOVeL02X/2hl6o1WN
vedss8LmtynqUtAl8IEyhyP2KVeY8mF5S47F362IcknNwf2moXyhNRV4MFsDfC6qEkjFw2wXLa62
cyQ1SJvljqChuJjW3NMsxZ96fUV1YJRepV8f/2JrTBCq90uF6A6Ws49PwLMSHGr378kHEAi5KH36
VVI84aBf14AwbTukRMuWKj/F9aFT32gVGLFGOpreJHx1NJvsYFnovlkLkBHRKxX4116grY7kHJcg
syYxe+NS1h2/9TAJ7FaaUZvT5AwIdZFSApQqSdBAiBiubWHjlvNtABpTjqhmlr9FuxvaaqXa922b
LdXewVjhhiZ1/h4+WiHuKAonBQZjNpLEoGg0TXTwXkfh5bNjtX7tXhYiOiiPhF32+N0tm9aRaWD9
tR+XfCkrLwBBzx6GygmWwcgqR4cKIeJ5S2c3pMMv/Pz0RvidL1B+0HmgjXiAVgG0ow5guV+41a8v
fKgrtH4Lg3aY4EzmoL3l9Fnwt2FZihs44PEgNPLmYbVQ8KB9vjV8GqzqOcVw0HgiGw3NBeH1Ac8b
V97UJIwNTIdIOVHNrcqyPgrBxLwLLfhTZZJ2qkbhDRCF5CKNpXvV2UnfouunJIjWT3WLzlbbn5+f
limz3jkQ2CrXG3eDC0paxo00KcYG9Zfxuyhza3wfKm6vo9G4l4H28iHwBcZdgL8nZx7rD4Zw7/q0
u6r0W5EVtCNangVK06xkSixrp+My1GFROol0SyZ0q/nPsyfaDZSFzazXM1tH2h6Tz+4Lhh/MMArE
PxPm6SiNOA15V182mxTOc3P5FXfg1eZ9+2SN4PPNeCqlFxYFHtZUH+EEIfaTJ3rsnGUQ5DlDzNEz
Kd6LyCzvBMEP4LVlGxlgwfdzky6a69NwBulPilHtEZvsZfwqONoPaVCxjxsgxtQ2z/sn+PzvolBf
Ki+DRshwzNnUQHjl20FlEN9uHY1hrfb+VZ/7UDZ/pc99uWOgj1Nwja8nDhRe2aJyZv9iU39J7MgN
SprxuzLBdhrk3sXGo6j9Mp263qad+69WwyT9sbwQRy1pN8FVOXNESdoDXo7aOvVZsiaJMgiLVqMV
F9ZzDmP/H9UkxjOU7O2cUN/cRtPplVsFikiYNHcspfU7MEQsQfRHeblgPzmnHIETOp2kTlLjOrqY
gkwfLrVyEwUtvs3zHXHpaP/E4f8jEV2Ni6EZ4bSUUm1KdzzyGPTVrwr9zJIyvqB0ioH2GBckjrdf
GIz0S93HueozENyRbNvT0bNh01zf8/Y9mzc198byB+YmlbP0Q0FBqwuQYPd1xt+8ImNgezx8P0/r
xfTMc2gu4fk7xFW5u1mTHFxKzrOdYswisPo4hwsIdgTOCnVxL9XLlgqjEn/Wt2AkuNadouqyBQC9
UH6sVEkRpjue9nwb93yFN9mfS62QPozDs9aCw04UfB9x1iQFLzDadHRUStgQOgrriJE+O/z/4ms8
/Z5FKYi6n9ZL41QcteH2FcMUkGXrmC4htB7SGLMogw6pRp3yba/EwliBoz4vW/mPY1uFHByLkRCs
aVOONjb/DPsGLOzJmxjjLhHRd35JxQYwhnj1dD70mtUKOGd6/N8I0AUBVSFGg6538fO/+90k6Uoi
FVytBPsep51cEA9f0AENHCkqtGzW+29t2GBW9AxmaIOm8FaQSy5Y6+aCb7baBnSiZo1Rkhh9FH8X
2EA6SLqly50bI9yLpO8eQJh4qtPogyLpy0qNUemnKxrh1y1BabYlKF/G4c0JEwEn6qu+lA5FkF+y
4ylUadLrB0mFuJFd1r8Cu8x9GS/OJtbVXBOMrvtbZKkSBTvihhC8aWDsKKWAaz+i9Ht71GWHkdJC
mvDPMjPBllZjngMrRPJpPi8+R00HhRo6PQhRJUDIE1frY3u0Mwibpnp45Ox6RXqnbTpMoIA6gkMF
157CkcA+14041KcVRcXgyI32TiPLwxgeBjfcjf1Y2nJ+Br9CVC78pKaqeV4ULNLlAGQEkCKiJwoT
5WiUcinqIrtvVzalLUiHxQw8VeUqurxo8k/KSJF5R0mOFI+6nJizOU3qcmg/EvkauUm62n7hWNJx
J65ifUAQkjBs4FFK5WuYNJ9EKE1vWUzH4efxt5dDuXORk0zZmDspOesjWPywlMAw1yXvsGvwhVZo
pPGrG9eUmAMJYSpOssH2yHMubuC2lFZZZl//JQxikJHbolaSFzmEr+Sq5CsqVG9tdsVyBkpWPNxR
l1oHURIYf59XQswxh30ESipZ4frqoBo2+HvLxA1jLlWy4amhuKba0Aobne1mRNsZIfnFFLzjbdrV
woqHZDfDBwC285hMpz5eQu2CYfCPrDHRA8zdxvjgb0iiRIZ20/F0GgSvjh2iDjYzPp4sQltTE3p0
nksBdNdP2dtD6ucwpgQo5hyBAezJGjdWl+JrfRZokFQhl7I6BITu/uABm+waAJQHZvQXewzXdg/m
0+OSZUL9GkeA2i8vx0RLBRWeqxmHS1NBa2/EdcAjmgTZcmitVUYmG+JIKmuGC+Z7dplSf/14ddm8
ZV9KqKp7n2juktaIOls0dq7vVy5FD9Og72dSnbSlTu9SpwcHdlJs4fAkAzjw3NLHNQgNTqRYrmQL
CjrQyMpAcp63ruzVAX7LzTUWu6rEy3aQyF0SKkdPApLYjhv1Idfh7KM/x7nPUk4DO8Kn1OWMy8la
IkKnZYhz4k1K2geiiQvWhmFdyXhh4Q0g81ylnvSdiMHBl5+smcE9O11e8R/6NHOecDqFrYFtvOBH
9CaotOr1zcpACwxsJX+Kqg/HKCR3mc/eLwbMSy1ZOcb4IbUEZa2uohJyizlns+TtWSi7aqtIKcVz
h1p+tm54yglRV8Mih8I2wXFq04p6+dNQcxk5SjTS3kqFEf1aaNUvjuLeglz1f3cgBMIeGZdYmQUv
t5wKmU/mr3Vk7TL9ioHwYz+9mznp0qWHUv/mrCRJJM+Xo4D/S0quLhrcchepgQaBhu+tHWUC3zcN
RTWxxmdsoHjewiK1h2fz1TuWyT/JEFaOtu0GFUK3tLYuTjvCdv3qVtuAyVDuNT9VztAkgojHDuxW
9taOnZelu1c7UW71qy3fJ1oDZbWyubaEmp7aySehWRiQRuJMn1GcG7MR/LAn/CO0lan5h6UiEXGW
94Db4AZwkT0IoDk0AfbdgJDG3WfEPsVEllCmkoNGdRe84PJRkdS2zkQ8nC2MtAaUICWjWtluaD93
F82ZipGha30DhxZCyu/SarkEb4IHG/hkpRehtsI7BGnefXyAD6dEkE8sqA3UzstVBoeZRZXTfOJ+
Nq6U/XxouWu8U/lDJrIHIMImNPWVGzrqYqCm75EjBwsOMtuMJAG3Aa6o44RMnSeSrYu029zMkE36
OVWhOB06uveX71lDI+mOeoMdeyf1FKOtpYTnKIEEF4+JuvC9No4gWkrpdnDaKNI1AQaxeQ9RDS66
mmF9cR9jSFgmOXjc786ZoCg0zwBOiUK497GrIRc6UmHX3rGVFmQpicq3BEcJon/4BnWJiAnmfBge
8BvxK2V6/TiNTerOVJDGxNls5AxXWVlCj0lZZ5tz1rdnjYVsOxH5gs8NI72LVmGHAW6xPAmJsNoc
AhxrBc/wWZqPqnrQAUiPSrLRCB7Wg1ww6DbGYVn1mw7Pn213nQZggfKcFBXav8oGEQe7ENd+CgvJ
oYTX34qyY3AvHAoVQlF0u3D97NJbqUNkWW1aXBe/euyXJ9Q9JRHs9j7hhNzX4QE4qNK813I65LwR
GMx7EAxUc3P+U/3Uv4kQvujPkTowDgNxhqJbLgPoTdu4iHXpYI05ulPK8SqQoil4bNmtSMxmxich
0Ksser7/BMorbkaP3JzNxjZhCp9mBZ1IYdBZ2NbIDyITijPlBrsUdgFyNeg6a9dh5zSF3WbnPg5v
tTGxPTqaNsIbW3OGDbZzb5FMWzb7RVxqD+Gjv9n2nuShjyisUhqVTIZdDbKgM74hQB/iGN1Z65yx
c7tZUwi3Fo/KSEJVMdOX1EzpFoAb9XMjM9vyMyiK2lOm8ZAoANf90ZExYRYLCQroysA5PCkUmpcO
Iw0CDlQYjQKv8qj8ttrU2XiNHR+jiNGvvs46TxWZRuvj2ulHJsxrOBgz56cL5h6cLVb+py/gV37Q
j/TqmR6rkHBlE1nvNgtAf89MOUOPpesbRrRY9O1jgeDuRHQ/IivSKwmF1dDJQdTcQUGOGgrelVwr
G2jGAtryv3eOtJlnLofyXgSkuCZ6Ulcw7W5JXdT6QDmfMrjuXY5CayuqQxoBnzxMtlIi5c6Z6goi
fSk3O/14FNEEHjmFfYHbDCZRyU8BkM2vjVXfA7rm3MjhXydysQtBMbCyhWFrHoAQiI2Eio4752Th
tiutKMSQeJsRE/8cSkcd7qjLtVhnRDSA1MVyjovc3Oh+7VgyX4k6vv1sXxNk4cbVoK2PihZC3/lw
N0x9ndspC8Nt0/UeeIot4PeuLi+gee8gGTx6zyzPEU2T4QgIwUqjJkwSYzvNoqjBIYofFnFIe9J/
DH7CmFZkDS5r8zeLVdmMsScMdLyuzbNvr68veILQ3VEK06FRSBa9Mm5F6egJHEm+rtfIN5mBE5bE
k9VncGrm/ejoJmvvc4WMKPZo7ZkR6SP98vlyWk2SkFkpECy8YzGH87YfYKBDSnIV8yhBOxNzmell
sP43sWXUsvTm4frY3Nqr+9kzRCA0I29uUMOVqabvoAEPINpXaT4u5+BLC98WYZerfGJuBru0jsEE
esbKHzQLKtTF4aBVc4X4FcP2+VAwR+vOrPlS175CaouC9PyXHtpSHCcYfXWHFPNVRwcwdHRmZ8kP
YXO1qjGS736Y9oYfSHmVAotesfiIvXJ83pRBiG2MYDrVivsDe53Lo4NbCCnYT5uNroMMY4MBaS+Q
fEdyNo0vftsjQgNJiXrCMccpBPvDrJ3pwCH6pGANwdn6urHiCJeeBZ9pF94jbFewRs0T4mMHbHDP
1DppEUrLKyP9dhaF0e3lK2YFeBfh8yxrCU+nBOb9nz1UkNdNXdUV17xztcUjHpy+Q3PEwT7XMZTh
IbME12DIOVFpkqg3JJWYgSgjdthszibeFbrCiHO/I60FQdikqvHW1mxob0K63maSZ1GADwGoNOTT
vUfw9IMe5p7MIr3hso+yc3V0tGOeknBy+6lFgWPKefMx/PMB+JfvcMPHE+4CWCV0O/9CB+lNwQf3
+UhAf6nsl9A15TEuWZMR56a5RAcoL83KqC250kFkTIxWLLEQRO1FpLtVIAjiknteGYcUkTv54eP8
v/QQYj6qgZBg8bL/D1dVJev+29vkyai5JYefhNdjrF1ezbUDtJzyw+WKXoJ5n4O8L0/ynFcGsoBn
8jBwU99ltCyWArSL2Jc6EteXvSTfslfF7CGlYoV+fSBDmwGoRAslpF2V9qLgtMNRK5GXDk8csCPQ
cUDr+uiwC24CczLt0M1lqYxUrnFuWK2mJKpQLaC+8t3PqDZYIvL4C7K+mL+Lq0dHBWVllcHITYDS
EW1rESZnOp5//B79iwFaAsm0xYM4U2brz4berIHiyf9X77OCjgoeKW1aiKYerRNeglGjtRg3E2cr
d/qsjoClLGKqR27VFqlE0oQfuG8vCuzMGJWrVyD+7maKfBxt5Q9Iv3AwjUkRsQ7AR68UG45lasDY
X/eq0ym8PQu60sbRmJl5Jwp7UxeyiA1uCSV7gLwpqsQyw5gVWQtGZikq+uNAGxuaGZ0I9xchNR6E
EXsHICY/9ZJosuJQbQTFw5d0KNpTylstRQoTRuwiqSl/5t3iqczsd/GmPEqcnVH+CZGw6Tu/CbGc
y+ag641ZCeeuJdBq1/puIZXco2TXu2KPU9xZsSv1QsyclBE0TwawMiwyxTDH29X4Ao0r/dTnHWdU
VFyBYOS8Sr4gUEbqoOwt/6PKNEq7E/H28fjL1Q5qAgoLr7hCgPFlLi9Be74mW803OS9KBKmWl+Wr
jhgNYvccNGohOuhaPZeaQFayu1RQ7++NZHwrV1us4KTbGBPYUIJTMun1xG1/+Su/Ib5WX4Ov7GXc
Dhx13tWG/cOfawvYfgNxSUXy3rMfMP7+G5egJEHCwbGSktJImyKSufa50nHFf9aoF/Hllf0bnTby
6mE3Z/iJGDI9b+UwLB/AUufTxrfqX1yyitX+jhMed/uMWTmPIY6aNTIkoTP3ldIXmE1K82rD7Cx+
GZHCWdxLlSA92ChDCDsG2yKGbjehTyDUKMqo5SmFTgnYYck5xX2kioMun2WBb4sWUsbciWYEQ7x0
obTX2ks6gqgwfoPnZibbOfQTcmTOqwqPUrkJV0GqI4kyq6BMuD5hQaxbWT3j0G8k/t6vtCmJngmM
MITBsK0ojs3rhXl3JRDH42fcOTVbg8Qw2VK6fcfZwbo99RA91kTPQJjHxXn+qV6So8s748wjhgaq
vMd8n7SV36J1a3Ti5+Lwn6XUtDKoN2SN0J0ovGktCd/W2iyicq6zF3p7RbJHFE9K0To6LdFsiCRP
XUGRReBo3mZ4SMgIHa+C/Oo1sEk+EW9YCqzrhhGq9p3HuhGi3Mevb7nlVpT3nMzv2ImuxYGuX/VF
+X9IP00ZRc9gxfXvX9fAQ73y39bVctwZF8XHmtLpgaB9b8/5BO7kYEYweuvxOOJmVz7zBJsqV7i9
irYgdpIM5s5Uytserq71IMt/vT0nTIKQXDh58ebR7OSt+xOhnFGs1Cu5Blq5/LSpllSdDLdiysMx
R8pgEn9dtVWMraOx9vnguKKN4D3YCVMgYVPcs6+cqvhVTnYRyEP9XX9sRVF4/r9061GjqUD/JvWU
WbKilujxv96Nia/aE/pzjfXsXEkrxAk+A2aZICU7HoIixO7bin0aCFBiAue74xEw0HK33QJnDvG/
MPTYHCiPXgEUWzY8BOcyodqW0iYMGUNwN+uotKj3V13XKhi5aFvVCt6dUW8l7hnQ32cn+sVrEBDP
/k39JMZtJUh/GK09x17JKDG2BRJIBRZwQNV0XHWzlO/7k1XaPel5W0QE97Sm/Utr64tP5qurN06W
1VBgUX+73MVBmYWWXDMAO6yU4Y1V9DRuRWNAToufM1VFsxc6vFX89EqJNSJWYn3A2mutxjHqJ21O
NPEGqDw3oMvgnspW/TStl4HD1md4XOcGX3AKb9B+sz64bxhT6DmoFZrHZL2b0eHEd4ctBEEt7Zci
5uy3IAESy3EAA85XBGWH/2NhpMhyO+pX0HeAEayrFiRWN9WCgDRLUe1ghJl0QBUY5dzbzdtgDUbo
DgCbrPwuMx6y17IKHrVTwmFRWotlc7LvbZWjQTp2x4odQWTXUlFkZ+N0WFRINDXSSs+kZa8d6iC8
ERFrYoFjNg38XQTBMmX5N/rBEPBIfzTrAQxHdig569X3yhcPfIe4s0cnFyKDHxCOTJL38QePA6Bq
gj9KM+qa0tOLW4azirlh2uf5gc7khfcRQECpjsBVI6wY3vKKBPrXSf/ShyqiifDKWS8YokcfQmo8
hAQjbKBqKAb3iOFCHbE7dxRMsMdTcsvbDqLaLkK00QOzg9LEBdjqz96wab0N4PHA/zeo6OUMqbfl
Nw3uf4qKUm6da5f5NsXmy4k6MJKdbJMxQE0jelSTxzt1d3bROeyeGjDtNL/2yxvdFWRMd8Tj5bqa
N+znzYJYFSPpJcGxvhAW4osQZC263J7aCNimkX7VMqYWjhDsI3zwTjmaEK5xTdG1siVK/m7t/hxi
LWkGyQyDF1sGZgt9Dw1g3hv/Pesj7hONA0XKbyjV6cBFsP3jEoUjrUy+hGMXw2kR/HCj8DudiEN0
GeltPIL4SPsP9svsPAmC6+cef7sFD0mdoLxwFbvj/PsAIf2L4yMUsmAl/xUeGKuwkiXlopw2ntyp
cL9oWK7OEQrWv5cht2HOEANKFmXsWb73+KthORaBTe/FnPx9AyMa5Qe4ZraupL2OoPRSUm3GxAur
30A+GqXCMV6e7ePR/ZBKCkHBxNrjwQg9mm0Ui6lNA3oNwnbHjFgUpK7QhLO2SDudrtMP7llzr0oL
/EzqYhD5Cj0w8NR9p1lP6nqp41IumzR5mn8Y26T2aGJSCsfZNpkPyLv68dKcXzDjU2cP3x6f4Fnr
SJ5C86mi7KnrVMy2wRY8vKKGDH64WK+VFaK0WP7pTk/oOVEBka88Guj5dY3JontNedKs2t4zOQXU
aL32ndYQKyEjgXfZ693HVUld9sHIiGE5//jQ4GJu8HzUbyQcP8LyyGwOb0x1Cj6WmV+mTtlDUnqQ
0WXfwhaSSR7b++arYMw3VHtXQ7j9Y86kGkio2E/4pPH2tQUSwUTL7dGwjTUa3TClKKGn+/HQX8Nm
GTMH7AWOHtKXZulimsN8uhQ9muOcylD5iVAfCVqQxoCPAe8UkMtYRxCID3+xr9gjBWR6+JH0fdgh
uX+FHbICjUEiFDoCcMpn0dh2a2tRf4vEm2PiUz6VckcbvgZinKp4A5/QYAbq7dgKqMCeGyNUt2DB
UoS6QoMrrTvW3smVWtz3NpfQycLspajmMJmzsEwF9lQwydhct1RZnOOHc+Ex2JaSHjbVujWh5Sgb
4f7DeDJDFctVSR47xZ/sa0bcf9nUv9b56A2K5QRhOSOzAWKmSG3GFzN51YuBRXg7n6pp5LG4TIAl
DV4kGHxZWzhi4u8OjghlkV3kIMrujR2XmH2lxJ92Tw2mtp5xTpCFv12c21f9BYO7h6k2aRynW1wd
cdn2dKyBbMvEko5ZdYaCfb/xpsfGjG6D7wwcj0BUKiUwsvDFTA7oo9zB3a8RJag7grgf5DjyqHhY
ZYG20c6gR26HZ9K41u9eBzcoHn7VY008OuO8LUuSVT4eP19MQVDikj14gdhabfJJrBZ11aJlWptB
JDnBQfhQimWwTgc40cVY9B6EkTsRY1hR0mk3OMH4qb/cN8pQt/OVX9FWUkaVWw7vknik4MKzHydm
NHMu9LnhptxaBbdxqo/IOvRh+heWxlgRJ1Y/WiUfH3XkTCGka1ht70/nAT2Iofg9JsM5nNgapIJy
SrZlOtHyQB6rOeNkkRXFA9Pn1y/J2M4BvXn7jxNR1T5w4AP3CnasL2wfu7u1Vh3sIgC6PjR6DwrS
iYFr259XMWsCqUwytbheSVuSFba+JgKqzQn5PYlGKs/fp2vIW22Dbv748uF/lX9ZD29noi+Y2Uh6
o32RpgpdphtQcOORXkVA5Yy1GRpsfDNAmxg2u8DmZbhNElwDM/4MLYO0UzGp7KBUgvsBHhHenZQz
IVCqbckwj8eJJWAKAxEo7+Ft5L5T0+orZlvRktkWVQv7z6Kdl3Jun2Fa3gdAY3SP4IQTTiPimj+r
E6tdJambXhXA/cea9NB7jBapu5g8xUfx4Ctl23y0jPt6dz+YxC7H2vgIN0f82WRlMBqm2cKHIyeG
cFHsfy0ImE4HKmAqWgaDFiQZb0yCMoibcv8Ci4S5n4h7PLSJ1zEwiPa+F6uJqTJ76jszjlAvXbuq
XQsfeVM8aL1WYE10Q5goYA84LFK5nHOUvm28u4aYmD+JI/qnSzb3Ng/FKzQO+1QXeqgaliWJfL4e
rM/eslaOwGHtQ3/nxe/lODYZ+NBVDMSL+Kr8oCem8GXwyvZepuSvt3CBDKJob5wa3ahQ8yGrX8IQ
VOTT1PhP4/vgLMlmz+893fWIfWn986Y1pFZ60lMmUBPgFiGGLC9GnKrXAnfkCaG3apxvRzZiUFXv
HjI1rfxe/nUXLEWhxvqaJSR/qj6X8xprdtWjknM2J9stRI+vEhlH22zKwwwu7k20ASnG4ZYqSUYk
OlP8CzSTID21jl0HvIW0oh71palSipNVw8cSFDdZUQM24GgEc3qlcWgrQdgyyxrdWEwZ0/Czwwz7
xhpOCzO4FKE0clJxWpDO6SLHlL/FulmUcYdpCXlevTZSR+THuy3DcvC1vNO47pslzg7vpAKSL4It
1pC4UVQhzZpYKIetOXF/rhzdA/pkan/oUw/saxu8rrKJKqrN04HMYMaHfQCqAC8W6DN9yX3rmSLv
oIPWpqZhis4hnyB2ECDDB8MmuH9ZJPhbg95iOp2G+kERcN13wveb481BkyTZoIjXQnHhFsn4c4ez
L9j3OIm/w0Nn45b4f4MMUE+bXbAECI9JNLLaoWnNyQ1GLQyg7ssGnU1hSXNRAW/acnmnuMZ3T9R9
BjRFEqjlNAZVi7x1kp5dlSimptJZMscIMn4zWVMbrry0+DMbbw00Psh6D7f/xAXYYjeLPn/KhFKh
5I3OaOszyHVpBpHrOp5POOLZuflrZEpmB24IEd4OehT49WLlkBt/YlQ5VqKLCXS4UHiSl64Je58V
cAK8W/7dp4/GsIyrWhkihgnvRBqQdnPLmE8OyCBMdedXHn+R+mGUa2uWIbaEUR+C9YRuutuS1+DY
c9gi1qiHyIb/IZ7jjy1e7UKOd8nVdyDhxXfRDnQRIlf+ruC6d4TVLiX3K0qocuhSK0PLP+G1W9zb
JHtJrzTEtv4nDi4gAMOQbS3r4IL1ic8lT64tFGhFO5otNNi49fKY24NivZ1+8qXoYi1o4BI48+Xx
vFjJRnuxTus1mvarM7f+chfVNSddjnqpUubUw2ezCj8s68BOC9zZXs5iRv/PxCtFLMQaoBSe7+2R
esSKiBICJAMRkxkox09belqSWly1BpiDN6cxZ0zhhXAGANz4Pwx9dNeqC2jEJ1hhvFYfrIcOvjLM
+S79NtPmdqegUwi69Gtuk3+oGL8iCXkawuKLLSCVzIehqzOOLjTQR2L9msSWLdFpRPSuA+oAvwcc
ooHyxqtuKnE5hCJgiHggLEhLZ2ucEXF9OnntSjnn1g9oVAYJnzG11sRSdV8poToK/uGlHQD09V7y
xqjutJQlUDjiTUw4H/eAYtZIeFzNAs2b8fwo+U2IosdptYzY/BakOBfhIRt3DGdcPuASEWLgSB/r
k2pLnx/JyBeWQoxPXTSSXjsf86072flRZg5Gn5QUZ/1rwiu0b8Ee50DO+zvftkRKDLAjrSR70OqE
BksdwYMNB+r1OvGdNMEnofNcfLFAE5yOiNAPyTxgt326+lSik8XD1k9iHrufHpo5XmamSPku4lHL
8f1su8VrdOC0dZBsBc8D7/PRcl1MBHGOqTRJmbOLqNe1EHgzNYCfecEOtXYQmCHVXK/aLiDKgGmC
iYhxtTYm5Tj+iPTca31l6u3rwd6/UhgVDBu9QASGZEOf7D2ql8Z/sr0zsRPReBZh4BVBNtN0x26S
xucGoiT4AX0xpICBzHyj4Klm8FxQzAip00EQa7HHLShhxFSXH7CLss0DmTguXlVkHcoxOdQzIHQ6
oT42h5vXLJgvac2ZkQMD8/nz2e22sxdS0YzdLFE/6hj0ZvNmPWmk0XR/sl1LGuJB8kGM4iBOhkBt
pH03dTdyE8NBU6j9Y//6B9yPAO7vxmoJ8Eu3hkrilbHCEJsrYpjfvdVEbPSfShMJoxO1DQTFPUwo
PBOYtvee08x5C8DH16gSELo7iTB+9OBstHQFkA1T6kCnaNuaksoiQ66Zh3ikJlmFj8J05MfXFX34
TPeYf5Fj3Xwe3T5xreTIT1lQ8bKo/VY3RSq3mJc5oG213ysFSYzb3B+BHM67Za20X875V+VU01Hv
sA8dghrGmqGGbSwN7oiYBbFOfpl8nkUctBSyN8f3kGe2LYipIEN4c168tsDDoPkmr/3DTEUouOtX
axKoQnk3ND9u4B+dI7aHhitBoboFN+BY2kQpbNLMHYcYEC66mzL0P1+bi6yVDtqm0pdT7gRi3lws
DDHD96krZ9XRKm1Ut8mydCDGftMegMQI6tI06LkggxpYGu+ll0vXh2jB/euLPcRO4dv2RVK+7vup
1cul0z0awRu4zmnmEGJ/W31Y4AfGUA6RCYqWv0wxJMQbr2+d1wZ/PHO03UuxOKceUGguQD6hFbuI
IEfmQcbVPST3apigSGIhHXKKfvbQzUnemJFBR4uZtqf775mYMqL7WoGFh83DmMIMr4xHkifMSZg8
W1tuTe5s/3MVp8kP4JUOJktYJs0tS82wqTme2RlAIjeZnbBit9viTOKgPbq8oW/LU/nOFPuP+zkZ
nFHMLCMBjGbnFpQAZQi1b1vsKCaiHvw/MC3YhzFp/17+rWhZXXKJ4oHFIkm0Ioqh43Pe+6bzVKH3
Mi3MTorhaKDBvL8J4ORPpu3mcOS0rYyfNCM8a1kAEjqGwegtkysjVn9d6DCZDyyRKRT4BEjoS/as
5HyvUYp0DXXQ163WkYd0hRYZghLOs7DWjwdP1IwCj5zXqxl4nz0qINftPNUQJNCGVecUY5S88kxr
NiehgkqQTX36uRiP4iqGJPlc6i5Cs/0BiGRDc+nszBR7NGoDD/oepOSnfcPQSZfVYbD4UmRtktPF
yhwNUbeOWQ1IDvynAg1qtz2+rBgkyzHnyP8VITTuf0fMjNOR7OYWZ7auZKanWd0JnAdHlGAIDGsh
EiSroGraNy4vNBRDj8rAyKzdZA2YW5Ghfk7yGlEUvafh9y18Th+gmO0TGBrovaGNgPEM8Q0TW+Nu
odFCUH5WopOtGK4qpwNjmF8dGjDIE8sKoaXwv6G/l8/oa3hfGMQSRDPR07z8Ds24gbNrBQ9VieWl
6DHxjusSzSnuuU+c1lqyoE+rwubvJusZwCuw2xmefaaqqBKYs8/Q1GXVOzwgnA+pNxq/TX8GB/uT
QXlCEUnfhkZJsySOLTs7vGQ4QwhejxKobppkS98mngF/lz9/yRP2ZydNlgR5xCy4JkgYziBhW19x
JLyPsqpt2bLNY0GyFyv+iwKvRqVTzfygkWkqPzxUVZng+YwBdOCf6JiRBdEytbYrBE30PGD+t2ut
PongyZVHuJCBzeUoJ+MPGpSgB0MNXfsXE4IR9qn727nNbJNs/XF925QOdy+T8RGIl7KXNtv5qNbO
8nzgIcT64iWEmKABtTMehfa6bTfCeZa2jYm/L2noSATOJM8+WCngygzinet4dw0hgJDpFmtDqmek
igDQ85YWhIE4CTZoOX8HWAbra/VQZ0gJGgidd1RG6Gvp32SU7tEKI6IhcObrlzcRCjV+aOkZUUri
o4s1QszIUtFxKavfwFgFPhO1o/UcqT8BpEOEr6SJlgo0sYUupnYCjqtVlyYBWwGbsuw1NpPWLTJ9
UnjQ1bzlsnWNKXNOaDdET4jCdMfOH3NpWYsBqXYZjegVHz5QfIRgNTStvFnJqbQGJ1JVnFoTrL9a
40x7j7IwO1RcGJns+dPToMdDA3UqLZ2L0UHtwY2jxwUZlxpVPUhI2i8yLggJVmcRq6PrI/VhpKU0
nOJ8IaxkRqMN8NZTb4QCZzBqDH7ULIxskucsbLr3qjXFRu8lJgaVfVXE6H3/SxAwoEs6ZcEJuiKf
czrlvb9wBUsGupWJclvV3mq+ok1qJDpDXzL/A6Uoew6EhSFu//99k8l8BiuhoGkRKY2t+9ubzfm6
/QcZdPKA/qnL00nsE9pFsEONXSalyJ4kG16b4rtTE60B/mAWXSqNJ517nECDRj+bwkwjOY1wiKLG
Xm0P8wb8anCKwHlZfgWDKNEdqdkHs2wn5u5Lg65wLWxLWctg49hmkDvoHo4vZ1xmyNCdDdVpzJQk
S0ohL4OZ0tWi7Yhz8L+TLrgRNk1zm/gm3ev2aVWoHfQCOKpL7FRLdO8YjPBRQ5H6j6Vzv+XDyI/t
wql+lnKmGGxqHZ0BgZEaSy4wqbIPsqDjV+bzrBkLDXJRoY9mqiL0gXUyWj35sC65ONARk6AnMxQP
DiC36LqUYi66U5WIR/om4ifmhLuCIpYbPtAGHWPtRmhW3zHC4mQaLJ3BpWsk4eaeUMG1WVJ1bxFA
2hXCBAa3q0HtlrHs6WzvrX4POMA5BIxyNU5oIQ777HSYzwPf6UT4JWlggLYKS8EFEc8kN8tFVZnY
yr0wBIzsMuAgl++136FJTCJ2qAlnLLSByh40pka7DX9FGCE35Rtrk9WzZjlJ9zQSI49kPTxjV73K
W5k0R2DVA9QLdof2L9MnnqJyRHd1M0lDpwV9BIGCHNKSk3op2XPpYesGi8ypcAd+GoUBoouOCCgJ
ALRgBfMWrvUPqzT1RIIqm1EW+aJU3NQdAaIquU4+OzI5AISan92pjgRInErXtI/pYmFFVoGe3RUj
UvjBrrc+LpqB2eqh1qSzDqRg0kmL/TerggmdHVaMqCjM9hbgaSBcHbQWyy0UU/Ep+2zVBq1BMP17
2Oi4e7YjdntU6nG1s6fdcHZGow9Z7qsU+57qC10pkFnyc7ndK5XeWjqH0qNgsxjbkgiJzR73ntSC
6P6lqzdfyOQV/ssCwdNnEgyI2SQGonuWpugS9QE0X7BHzJPRrsfDqGaRx1RW7DSaYqQ4xhGmiZwT
4vPyG2ddSwPRDFdKx8HleE6C0kBGJ5JYtg6aZZWTjv/LHTN9FI/migB5umyXmmxpKr4+uxOrl6iu
zAmkDhT0LTBx6EOnUTRUYVYF+lazpUbWWbqcOfqrKkHjjaUxW9zwXww98zkH/VgZKYCsnYBAYu3m
elNhdpzI/FTCicWJZyORgKIl/fczzRf/Kez6DDuIe5AS8jwnTDxwVdaYULrh6fYogGUQ6c/LKPae
9nrD0nGofKuN2AbQbedZWFJO9w3VyO+Wf/RclyqLWjUAXAQea9krFhYIItfi/Nl1KTPcXaLIEaUY
ozFUV0qrchPJjkA3oh4HdIaYX6b5Z6Ah6q2HGxWwfSFh8EV9xaW8wYvowvV4ehEy4XjKMw6u3Yk4
JiishVpW6fLU2+pIvWtXFgKc+PRFEEhYg/zwOQ+5UQsZFyQBlBi+vy2yV4jr6yvCPH6Jo9JpRcyv
2B+hWJn5cM998bphZbbVpFg2j1oBEpWE1gbI/eCaaCmbjpTJ5FaBvdS55ZOfxtCSFXkHOUlzH6SO
2PQ/R7uyl7yuWkiwuPsOZLRKhKCFwA/9wEU8LZOzB/yD0Nfxi9zbOdbg6T+7tMHSZ2YLWnOl6xCM
uTbv+L8jfrXrkePCyMTE9yuBF50hPNG3JUxUNSyJ2PzTIYB2t+tnPcAbzqG0Zkz6mvkwI7MNlyB4
TPn+hTEME9pvkIEq3HkpJhvBWuHwdJ6OpBHjf7ndQ3xWyEMPvZpfZOra4AZrGq4VEybob/FHQBtr
laaGzzQ1GcJqprau9B/kUxjHh5JkM/Hl8Via2PI8DwyyiP0/QtO34+wbtfd1H1G65yv+8w/n6P6f
6JMM+zdLqnlV/VqZUG6FDGe72LRvjJO8psvWdcCM5DNsNFs++m0/TTvbeq/gJ6vmdWj+KaOm8B0L
1h1qbq7Pprq1LxoZIiOPl0io5nInFSRRsaU2SmTHyvioWmtMG7eiIsfOsbn82Oesr1/gd3EOIten
XJKhXYCcHbDU2e4vPznvXFjz6FMQFlwnGcr1G4Ej/CN2NSQQwBcbAxyuKMys0ZAcSrqdIy/tbCUK
tXGa2k3A1qJEVJ+k/i2tLNFx//vdexYwe7x0GzOnJOgtpybTOzN2OQsi15CPtIpidJoI5XRPZ2xE
OmNe2cxYdouqUbztnx0BJJhNkJSst1Vfua+ts1sSU1tp+cyn273rcHkWVIrhqx42VwRJmot0A5Ls
+0T3Y8kpYcvGK3Z/tbozO8drwSUc0xgQ1loRp+b0JF7EbK2flEk4pqQTqNIc6+wq1arhhl2SlHnI
azaTO2Yazyi0ZRW83e76XiVs0CI1XL20fq16vh/kuDJPfKCU07742UamfnxV5ElfSk3iGIrfdNP0
PlWpUQc5Itzk1ZTsDZgd+cw+RczdhuxprSsNWbiQclSpqnNSib5ntWiKd+24PAbwT+3cZkdZ74S9
BRI0/SXx6IFgEemdANvIX1TrwCrB49iu28PJFlWzugI5kOQRJeJR2kgQbOallAqL2id5j1DDr9nP
OqXW6GDaFkK59ntE2k8KSLrffKD7XJ/D1AYIXzfHkzyfHMg0yPgsLW/1FOM1A5gZCNzRT9jSS7/w
JDoTfexcMeC7SKW/vktMmWvdWKNvHhf7WqPMgI8ZWZdEQSNnBbnArN+IpT6oKLqug/Q7neazImc8
r1EWf1p902UH4JjHwmd7L3QWaKaR1sE/u+Uy3jtJAE/zIi8b3BxfhSo4PNi5PZ0e+LK1vQIGCfHp
8bxYkxx7xTjFuJstH2WTtJj3V4xpnI/JmPSXZhLYtQN6CPwaf+z4++4k2sMGn0oXU48SAgW6HQZS
Ex19oROA0Jc+SN2C4p4IzZasJkfv3X+oG6uAtO3czO1jyyYIIfh+XgsiTjBG4KigBqv6n1ii60Q/
VJMjePwSiSX+Iqaa2s508Hn/kn8KEgWBGXxJpLpJzex7Za+xVEks9vctZuuwVpcnXdNlSyvLvz44
hPel/1YUpnmcrwuyDT5a/aXRRxPP9mdpe3JlfKxpc4DC7wjPDYr4yS2Q0bSbWBRjAr2gIfJGmZIL
gB7AdI326bbAFk+x3JsERpQmi0wwFsgQhvkjWEcnJUjiszZsHV80fNXZvwrDBBz3lflLpDGcAH4m
F8JVDqRX88DTd2poSTZTh3BXcTJ1HJrvW5eDTeniefOvGjLLCNo0fNzY9SW4n4lr/aDHdAcIUZll
TLF2UDwopamDKCeyiDFRQAjUfRX0msUDY9SfBYaixfQ5OBncaiKzvCXQ/K9UjudSbrNIZRlNSsgn
AyZOCsra8Loc0+10k4H5I6WhCwALBSwxK0a67wxfoomR591bN815hiYXFfC882eA+7NKJPk2Pr9y
ukrCn/jVkevxkYK+XYXt0CENg3sI8K3elbFU0XaD1B1+wm3MA5SPmilTU4YAWy6zMeUjJplpve5L
TjEfOlhOgfT5xEIW72vGQB6JQ2q8i4BVD6PGhOwZqdNAtaLvQBVjKoe1+8ia6tZ8DrnwdY6XRCKF
bT3sEvjogq9KLDpYTt/vVLTjs6UqBVTqWobJ+068atmCeScw9WJJIpKmHk4t4kb1EyVPxpCSTZ1/
dOijBWRXG9Q+WanRHyUp5JJxvRqH6Ixk7Va/FDWAosQ8XqkBfsvsewlQx0gfd0tsTbNFpXhcdRWb
ZNbqBphtP/HImG/c/Zysyxtug7Zm8DVr/j48TjQFFTNHu7OMhIjAfXnoqf/Yw0y71JviOzxxOiHC
P2WpxCElEQpxRsM7I93+MV9/DCJcUOl1YHBOWnNL6KFHBOCl4MpDy78sNe99tQd+HOaY4aSxKwQO
EaR7qBNxRMh4nkpEVq8jYw2h+pbBedw001wvgXMOoCCU34oRU4ILfXzdf6tBaWgRYKs+gu1AZn3f
mCY9Lr9I4T68t7lnrO45T79EHmh5erT4PuHTlueXFYVolbRawEE2Ln0gQGg53fG17HgEPqJlwQbu
fAplbENRvj0QRCmGp0E6tfAl6geU8FjcJvf3yifbJ5YYk5l1CZK18W6PzbrwUjtPHrGvA+MeKhcI
LtaaGjyYgTugf+rZX28nb93HdnXeQ7sgx2CHCMKPo4NdP7B7UhFFTLmEed/92hzAU6mr9Wrg+oRm
13i2l98RpxdrLLYIOUMur6ADwILJfCBgRjD9vYnBegTSvm9OXNUiL3BAITXBfFShaCbuzYakHMpc
oCXjSS+2Q+e8FOFGY8IhSGe/aQK8FAQrpXTrGDhvJYlvFRX11VLjZkXvNSTb7eXe9iZqZ2pimm3s
bnrDSTG+hu4JwuNMfSaTPe9Qy8qwdCx8lwX4QznR0zDCwJ6NEY8Bc4CDWRJ4J6dDkgD0jK9HvRMH
7hH0P9SGIvoCq9kkQXjDN0wt3u/8Ad/MbhfWRhlakA8afkGBJUrGR7U0BSUj0HYFndSZ1cqhwEqx
YQIqhXkUtVWtADqFIELL8KCCT5THiI07B2suXZIoPhzX0hdtymOxQ0EMD28whH4upOYDjpVgY5FB
bfeKuGcwK9Qz02klKrEVjTjJukG66eqsiu1jbF7pG1VGabSHhh6fDtS/AcE1nJ2Y+qm30R0JVNaB
miljl/UJclsKr5oMQ//x9yaZvrUkSBOJ5NYxPA5dMDirl163/wQrXbkkU7+DsDdW8g1Uwq0pk2Ek
WGBtFSmu1ZWLo4X3Wir4qG8NCXpgreC3XNRH9SN/OlUru5n0IsWdd5A5IWrl3wRCtfOJF4qef1Fq
OzCal5Xxy8wjTYIue0IO29KTPLS9jzGhJeDvtPM4OesXJAF63fZvOIOkKuLxm49dnQQhdbX40XjH
N0jVP73IQB9dMCS207x8zKMf8kQ9oRIIWdFsnrHue3U4EMKuqaQdr6H0iM8FSc+NVS60ZvWwdiIb
e7UrlyTKzwu3peXgA34+TP7wouEJ6u1hz/TCp2XArJaW2VVC8JWXxESC5pizX8+P+DoLpAYl1R+I
Cc7uJfWoEU96rKmFCOAOcsFsBs3mYIrhWxiOWIOwBh3Ybitrn5i7JixNhOQJdbfOrJcgJVGPT7S/
HR4L+DAf+S2C/tXTkdtXYsYshPmyPZqqwHXFCyEDHfa8vprYx6RDdkFYQ+cTog45Dh8uNUJVTtEI
zl4NiPOgQYCSDDGlHeqrrRhigP9rPg2ofDu8LKZxhBKcpweD7XjbscNV95p/aR08QDK50GQn4HT3
ghbkW2buK2YwvfwKmZZU9vc9KDye2SxyntCkPaIMuZslZfZd85yzqpn9zIxlBd4pPO4LTPa6SMVX
W2Y3CcA8H4iFeK35AZV1sL8A8qTRcpxFiSKD/ohL7DYaQlo1B//x5eKY7NHpAyGJkwSsEO8Y3djT
5fPL2RwHw8E79oCO8I+OvmjvfWx+yNjg9R6hJ7qcnAfCocIGsUIUHypvnZ2quajn+SYWPjDzYZtB
TdwaPqCS8qGgT9TH+DAJwbkHhrEIniw354e0gfYSN93ReM9FZgYes/BNwTJ3x4DfO2EZbFWfEaov
DifD+emxaahU6AC3hQiaAcdI1S76Q8s1cvP8GoEGfVmLZw1A2CjiGgzvLhoICcSHIMljTap9RHL4
QcN/o6aPBb6Kojg5ilnTd/CzKndisaQ4cxaOxQGXiz4ky2c/460WG6JQ2DOEBTaPwqmCIl5m4e5E
pkxEBAIzYa+Cs8KeZARnD+3cZdnUh5xGPtMzztP2FoSoSOUuKag4wD/jnlgFE5bBwgD8Ckekuiw4
E9K1PfkbD4qhpeqAnrLIt5s3uDgmylfFQGGJQSV4ia+FFIIYC7bQOd750ldnlaNP3m8/sVejiQul
nkQXaEHSkA7Vl+UnnMosxOUaklJa2RgAbBUM0DoEh5GSgwxCcjkI2HhRkEXJTs60QOqTDZNXaE1h
5rpy0Bnnf9PabFLHpJ2ktBdOEXtGn9hZsGcbrmDOjgU8OG5QxhDkBHgZQFLaGBguv78yHUL1Pdd4
6JJQsQqafhkVgamUA43BAACdDMT3Q6ksiYk/rf1WFCL8JaN4Y8fJ06wWNeD0ZZMuJyFmHChY0410
y85gcaSnzRj9+PejNTmPfvDt4rUSE862I49vry9cj0inWl8AZXQ+OXe51gPnE1dFmSBC32+KSgwG
NfrhzajBKV9BZInHcx/DHL10AQjPtbrBSdKwrd6jd23auUeks7q3IqN7UUlHIyYSxD8VRRGo1JAr
qCnPfDLxWsb7JteoNTQeX355hzo5UvltIGLUpl7ALXY73w0eyjxg9E1PY5RIlkMC5Ke62mM6aGFB
aASUYKQR66lz2jnOyuWmDzR1mHtLm0xkuQ8ux6/ZNZtDORqHVMQN3KSHf6lPMXE9A6+0K69uKELq
09FTJiS23mt+P0OkCM5ySl02V/aRnrXMFzLemrqCHsHWmrr0gWI47N58IR4tSwxcnPUcYxt9rWMR
eQQBu0DjKIIQRo2Ett8nLohAMYbA4OD1/oi/ZdUBHZOdt9qXxI6c/CXw4G0wfs87m9jPvzTCc2K1
Vot2u0YunzHun/PXNLjsZ9gcGlHmA3C6LIKBGF8lGw/Ao3ZP+kd+k5rjrgHwmSlmCmzxCsNwJ3cB
MhQ42dLA8UwrExIHq13JQh75cNeugUh0JU7CT2xUA6VokZ46uvzvUfZLGa2uzguk+OUJr+v3ypt3
Wz96kcd7fCRKxdGuEcXxfFDIWUhnEN7N7BfiqX1URP5L2iNc01y16BedQNqCtyXNSVURdH/UYrxf
JR2bld+TU+FNYnfczRsDeFhb61zWgdJCgwCaQraLO3DwWeVMJGU9cpLilfYjZS4pOo3VvFHJACMY
TR9a9XRwpmo6zOXWaWCNYGXkoeVuYreRNQJY2CxPDt6XGN0+FpSZTkkH7F9T7iWImGSpNkRmNupI
KLR+W6NS2QfUly9Sy8xwWsdosxAUp+XPdMDqJar8UZWSML62Sl8IMeYZ6+fbeBzLLptapOysapkD
NgZdpCukBAfyfenzmkcg2w+jwNbPTfA8mpNFDMLBjmX6uMxJGv8W70QlvFEXWTQev7JVOKXoNLZ2
K4KlTu2L5pRCBPWHf92g1IWR74NB0D6rJgamsNN1BeeyPsrnv5IELgJGs89I+EwnoMfNc3cIj4HN
G6UD1/acYseEqDVT9ePieVrcuulMHUsey5P7kI4WL9bI4wsdVjk21iCu6ynyDd4Y0indnC5ZcpSd
uari4VeRUyJdVAe1I+xD/iMpXPsnoK0DvkrITBhCg3k54/3i5OMWuEyIsUYwy0DEVd/OgBb4pzPU
Dob741PA0a3AJBN2Q1z954pVyJuS5Tn6CEf0QbBViI4NG0A8b1qn44lCqwOOZwYQ3deLlfDJ0+QC
ht3kE0d1VijiCceWOPNofIYGsHrdVLEbhZcbc2weXhiT1e2of2NqGlRBKRk7s/sUjMYK/oBRYSt7
AmiHapbb8KzD/+DJQ8TywvbQkN8myK96cEJBf+/TJNcJRhNs5R4CM+IlY1VKUaliAe00o2WYaf9d
ACqY5bGuiesAhzTE3MVjYIWdiKiFSdSgB9LZ9t/MEm95Qi8HuCf8ahYHVrW6OAlkohZhTOhj57AX
+d8JKc2jp2VbCyDuevJS7I481iE+4b3NpJCx32qrtZcN43BYbHH2ABOP6q+iPciC0wlxtJ5oj1cu
KtOM8fx9LR13VIOFm0H9II8FPBXZ++qslXkVbY/hPoNoQPmEXxU3TOwp7xR9Wr50tBTDdL1pU+j5
jjUe8lgrlDT85leI6So4hnqq/nx+ffdcTTzFaZnIiN6V4eYGtD4TKdHvS2P9lNGfAoXZYbx/ervc
4hfcKl+Dz95GH30N5uSniZgeB0Nv2Gi/5+Ed0qPyGEXW64Sgz2OZrthhpOASWFXIUyNKlhzW6U+h
X8J0Mf92Br01kRA+H28j10fGw8SC5RtFKoe2WryHEkVtFqGIBAelt6w5JlPidZoAkYzxxy3mFXLS
nARaO1DLbG2g0ITIsvHL/M3K653YM0ECjDikLMbezDsK4LLPy1rscbL2Dsouf9CToBzsAteHiMtB
TISoMFGdX47gKf8k+TES752X6BCHm8y4PCZ8uS+dIGZcGS791EN9iTn3sv3srewlSOyB1sxWc2xr
SNrNyM1fPMwdCd+PyyiusdyD+TcDRyyHu9eVDNit1IW6ACudu17xfKQhs3mtvc+L1kOLBBXUIpVo
Abb/EcVEBH4iqEiMiNijNRAJGaBWPNaBMb7icHtXkYPwNI1rlc4f6r0P1zbQr7V66PXilU2i49K0
/FhtZBJYbfyIYQ1u5a98ZZM4vmhjFq2rT5YFhst8J7JWhl0ZH6X7ZOyMgnXdGRfQEsblK8V23twR
XwmpUMazzBRe18T/Yadv2XoXHsdkP/2CYvEYkqy4zmk5lXQCVI2utloKfMWCi413sVzGDlTyYt9E
cd2UxFz3QkbheutiIPclxPZqf6d8gYb0wVwYGvS6CXbw/IxN58w5M3UkHCjEA+/ZwOWQvVsvrCJ9
7R48vs/PchMTGB0vJ0/26G9lPYHEQM+VH9F1Ngq0J1qeBggxmTxY0847CLE/P182Z2xJc9SPnTM1
Ms9DUIQja/wbuRk8MejxmniO9xKl8r+YNgkdswAoMFsbqokYO1OPZXqMG6Z5QbgT7RcuYZp9aqeF
FiiwK/lHdVPDGJgdwuX79PaZNMPLSZI5heHloH9MZqasHUoZQ8XLDDCgaMexSvNg76ZTjp/kXh/V
PN6EYp7jEBCjh9qh+EaNij2xna36iLQ2EVQxcARv96A+gYwdCxDa65qgVt/te92rr43AC05tSBAU
QHe9WmZrWF8Fc3CJkSimBZhBQIYSh+txI1UenNYy/H/DAsDDizP/aBud3gi/6+39CdV5HFprD84b
avjf2UBxBhMessxGTYdB9sOh1ejyl/fed+30467x9UTMeHS+b4qRjG4tyMW2zF/gQvekEpddHwM5
KPyXAK2gB8x4JyBV226v3iq7p/9Ziqc0N6EBeqOrSb53fGlF9WTTDZ0f9AnUlSId5kM6DuYUt10l
uM4y7SqOtEuxAHNJxdxddZsY+sgAWrHuDntAAruiz2r9hIV34B6FCc0YM5TT1a0eFZbJNs1L5qQl
21mBqCJlSkQIm01Ei60f5zZM0fjwZxVFhGw5xSrC9m5N1/tU0ebAg+3ZsrzrDizGM+7DMuzVrfkd
LZvgBO7y43PSpHkaQWTtW5olJmlcb9Ymue8XMZ01931E8f2W/FxZxNTTaC2N4jvGvnL+5FjyFNl0
SoE7Q6H00Ha/j3sU4Rtm4L4N20NFbffRHjg54RV8e3GWZAsq8jqC5rCMn4Jb0/gSert0pxtDT7GZ
HLiunQj+QUDSiLCUmDnuJkYvlnRcGfIbP8ik9flLvG2rXL9QrHnlSJKLZTNg2KHisom/5uT8SWDE
ErQBg4/cUeQ0v941sHJ+tQNTnXiqJTedQGBQjhAZmzNvuXpjX/tvkrs0/yWpMxb/G19CgSEoe+N2
MsKvQXrDqL/jC1BMa40hyyyj4/DTzHHzGnHkZT2NxVkEhSp6V91JRrCq5/E8qigsUBvkZ11LprL1
ZJxZEhvcUtogEzxPkXbmgLWy6NX7CUzeP/uxC9VG6M7OehHzuPFlvYfTpn4ua1vQcIMviSWrgLw2
FmrhxunbD/f8MFjbgXgpoKw02MmioTihw3mhSNa4dlZPnR7a/jTQKB5r3dYfsUxj7w577dESxmPq
zQwzPwif2T/97QiJ9Qjx8DbiEF7w1DifPkFthH6lAqc/2K7A6xGjuwc2P8DjeON/s8Pb7P/mJ2w5
Zhy3Maxgv0+HFXcyRRItxyhSlsUc60pObjPw5kezBh8+SSuIw6XTO3PYomvzuFsHT4O/49amFvMN
f7gUb0w+jXKpVemVOOJm9lGUX0RDVesg3tdCuqJCxapUT3tKeQL69pfhCbehkRukk1ViuPpKYnye
ZUo/RNPsn4kxBerizETYCMTPtii7Snm7Zo80Gv2gPRVVYOf3TrJK5ep4Z4zMBMPiAiCCgZ15+xwj
VIP+kAq54XCYIdxwLg1PwM+F/4p3GxrOrIdQC5D8x0hNJcy2gbRsvX/hjbjtK6SZD+ZyNWwqn0EC
bSy/m1CdeT9XrVtPdvz3dASnv4L9GI5PhkasTW4N4QmU3piekco+NlvvS49iNUMiqJJswIe425ex
45MAn/8T7bY/zYl57qCBCtcXHxqDNJJgE7IsJIptvNOjYfcBjt1IkKuFRZDAsWT5AwIr/D0ChlXn
073uChTdb79j66i0AcAcI50/+jGySdN5UA+trIaCOXH4PbZm/AgPu/BXN30GVkI/Q1blT3QCo+50
0sf6YggJZTFTnnUMeaNC9PcWgMb3fSYDIpqrl84hTQcrVD0xhPliLWlf5EE7fggv6MD6OsCmUNi7
ENVww99ef/bkJBYbYATyl29nR2en6yvr2vh5bFsSRj6cKF9T5pppZ3GPC0txvg28spge9uvSI5US
igXth7+eFb/RKaTGBy3eBCjDunpcmDd55c/fabSMqQD0LoGH5j7zyQ3FvC2pmY9zw8NiRA/IohuQ
tlvHUFcIPR6gV70qX4vw3DAUD/OclWNqX+aElO3CzjFsGpr8yiL+Ptojtr+D36OquEp+99WsmMtX
GwM1nXumEJgXr46/uiyxIwr23MMvzb5Ty7uQWFWf/rRON/yZ+OMsvXj2N1gExzFqvgx8iG2SGYht
fi4UtMChBF4PqglgE2zwZKcmMOaycZiCXmkY98+/MIwZoClS9mQZ4jrDCl7hufzX9tpJb8WaamqI
HTEjmghyVCw0/FZUdmWL/zNRxD23yZSXCAS/fhJd2/NdiqOr8iJFnbwTZ9wp1VJIXTQYOts/lCWp
Rqinxd/bW624aOD8fNHFbwkNhGr1q+TuvOmN3Rs074E7nuWuR+OZ7tyTC8vTHizSRKLQAUhUpSx9
42d6prZTd6SdyPXXSoL1awrKyQ7NV84dI8lXbNscpmJYHC1V2rN7wVjADVrOGk01QNAFjeoCs6kZ
NOZLy3+Gz2/VS3MaZljzTiz6rZe0/tB/VlICmkaijmQHAf7+KoxtP1z3tCtscgQJMHYzJR8qWCwE
P9z9/80AQCipQwIfDCoDyM07GEuwb8VtGjeYe5y6Y4kMO8rdVWXquwpXpupSctfNeHnISGqvh90U
FNIz+qDBSneLB1k3r0gPhJUdYp0l+LjfivAvkN5kN2fXMvJnCRMkHAq39okxIzqMZ9eWxu9+j0bV
7HhhrztWNScZU4zYBmWeFRiwLem0DK0NmLSbDRA2r7Bk2W8oGaefGahyntNipC489zET9avnkw3D
+qi2IlLR1xLkNIH39YzxDuIls7rLsW/Wgkr9fIZT+q4t3g0TefSF7b6wLjvcEL7+tOawKtzZ+Aks
/iTIQh00c83OiA0vV8uGK3xBEsGFFInETrGuSf1gw6PwDQ5gZFqNMivqjcfybkRP9bbilXNw9C+d
n0W38YVcV3MOw0KaCnTRlGU+llK0pFg6FtOA1yTxJTtquZKp3uu3K7BFrvpoyWkAc507gTuNjxfk
SwHjWg/vnwpMUnu7OjZzMDoZroP4GyBoCP+mUFFeaIp9bACKsfs1wfJr9rnVTsjRZRMWsbSK43L1
IYzrnoIRpCbBxqvmmlVmRdlknWkVVT1lrt5z7Hrv+yNAsCEq3bPNiuHlyT2haitANkr4o8PNP2tn
G7j34J8t3cL8pARnSyjbDjcRdxLhASndtU2/0RUBM9lfs4hKkxS3Ekyt8bCbAiXMhzj5MnY1+SFn
APnNdggcvDUurugaK7QRg55wEuK9W8mo75QPnAcSYKg7ZP50kQwvQrF3xH3GtZezbobk0dyqcBKm
9bhn+DJdMkrluyJ+0+Ix9GN/FsSO6pxqOQDf56djsXqqPPkiA3Qw2xKmMBnZYEly7tk2gMTcbD4C
gvTQ3qgaXN4U84HBzC0DgemrsMCo9r7i8SnnHmDMfS2hRcgmCqXA2PVW4KenPWkfBDv2JLvVXH3E
qLd255lOn4O0VbxzLftVMnKR4b/GQ+AFm7n0povj48BWwdeKoMIYpETnzfP1ljx9Jrli28lLRUCS
nVGsBjkop9PlmDL12WNsb9xCtFNi/DoHrilDjCvX2UeHYCFFNqOHtSRuODkk0YQMMzRYH/DtToOw
0i070hX8Bf2uwod88ECAuHlDMgO9hCyaZzVVQXRjVd5kWEjlRJAM3CsP78DBdKhuDgRLv20Hvq1+
eW9lJBNhLsm+l2VOIp+y6O4y1ITqUcqIkQIrf29Uul/GFmcoiqnAgEhKm/znLCFhKDD42wVNSRoe
KyZ24uTDhCs9Ks7vDyjmOS13BRBDbSQSQVVmfeSfIg2XCefXeJzewqOihkhhZslWKvBcO0rrbc2z
C/qU9CM3be4DNzmo0J0vRGK8UVU6JHIvuO55N9VcBPldwjpRfpW91qaVBGWU4NUMSkL8ZtjYQ8D+
k125Qw5BHyDKLQdZF1gjUSuZOgalM14ZHYmg4UQ9A7iLOSHwxnyGRnKKS1RihR/ymWAG6UKm72Tx
iq8LSGdu7GWBEcDStKTcJBV5JE8Wg+EtF/DLyjUgD0ZvI6TP9xmUKKCNl1fVvthjCScBYKuClb/8
nf7mm+RIy575hku1ikOwfSPiKYuiLTGV2HVCq+PCVDUwDWkUpQ7MH1FkPyIetpb3tIk/39BuVMxP
HLGdGVwYrT5P8nakv3Sfc9O8Za2jwvYLoHszxcE/jh0POSFkN/FEXglW27G1kjRSdxHD3gdy9s2Q
iGj9LGz33a2/R/Ec66fMRijAQ1LKxMs1gZhsvGKZii6GNqfhLZ+oFh3drRI568Ix7Eua4ewb55SI
pYuicvwlk2lRT8Xs+4J0fb8Qooq72qTdVlQiKMIv7SqnGYfqT+9WzhNQgnz2GDUbbsb/jhet4wVH
iZ/1x74F/YB4E/OFkdqkuwv8nWxz8ts+qQyUttWt4a5zwG8INo4lqDa6Eb86EP280wwKKk03Pqnz
h3llE5weohm2eQvXMjf7S5hJaVfXduVMAgQfHc0rVT4Z6f01hmwXaGqwfh5yQS+8ODKsn0rcBJdm
D68p99CPC776DAaQiN5+ZdcKB/pHJHkvhi20aODugq4ctH2a5eUs/ezU03YOAZ+6O4Al6kH7roU4
g0UTjj7/Wxi/KoXPuo/CR5e2ykP0HibpJd7sJA7NPRe1d0ObDdaFm7QH4f9iBNOSU51YGjE+FgGb
wxo6y/xbc52uqC1+c7+GPJfBsX/0TBej2Z/1XoxplG1+VrhSARJ5ylZ1/acsLfsD276wCW4ZI4lO
0pA/mWXGcEHSrh2iooifLL8py6eP71MeUAuARo6tlsLmtkdok9ey50cIp/UrjFbjnauqqqUPI7WD
azw34QSC88Qv4KSopxH3WC2VCCFJkaHxUh5K4ksfdEbDPbQVp85uL6UGzhPQvNNR9ScF0tpBGN6W
8YW21sEd26JjUKoAvuwweCitFrYav7+iAAyE4qKDafquJV+z8ZGUG2NrBbj+rEMZaPmNxAORNa6Y
F7E6+atVUgn+RJ9+Axu9xdaI/LVguD1BP3PufMO+MxAmSV1W5rTU9nYYf3Aar5YdBfFQYGvyzQZE
fgDHW4lbqhHyiKmZxb7YHo9qEylnLFNJTxg/XivYGslEYCiUwPh+gx2lwnckiJowQP/ejK6WGqqn
E+x5Mkz92ZBtAH8OQTo4aHkRc3Ez3eG0aSrn/OrmASxHZi57pgKcCPs5mB39/aLciQ7P8GrLGMyp
qDQkQSiL/0QObhK0D7cDzXbKA9LnM2Bi3AAo9Vul8rBRNCRzeXe4T+sQBOaKVXMaUa3eDG4LnGFb
nq0IFJYVF1fuRHAYLlMQDxUSEgHtdug1sy9QfrGuBq6iU5/js3nMVQ63gzra+WPm2isJ7zm/db7R
GjnFVM0NdFH1FbIomMMABAGEc9CdYOQiyR14A3G1QrUjNRlS3ywH5Ql84BtPdYzoXnEYljQB+uXA
5vcv+Yypm/qe17jlX5J9ipeF5oFuUUrIDDVQkolAYyz08b/Zs7yKxMhsW7PPO9Q5rXIePfX/3/sQ
HeTbaOMgeYEejg/BoKyUcYVN/e+361ogdu+a7pK5xBL+/bDDghwJpxH7EqTQPAR1651lWTBMFY6J
Nu5kwT3zwNWjeTK5S4xeK8AJOT0S3jZKvqCMC42f7vW31qotVidR+xO/gSGd2dO2kxk4lJx5LzK8
YkGwdltXOgSJazI613Bg0cdNpqoBekqEeYAC0pMZibzfLIxjCDWSmsOSApeNb5IGqk6sD1o42GI+
hjVGrNEDdqs/1ch2/BIxjVFx00bz+2eK/19SknQ/4UT7nrky/kNcYaACmrRsJYY6xESSESo1jjtX
Gb9NnDXtCNVCleEphK281/QQctUhpLv8osgvVOljM7ksKAnXSBEJML69aMiPnbjjax3wNI9Y+wbl
MpbekTvIQ/qW7Viia9yxgtyHf3DMtkKOAYFKwq698VeLVoth7pnDEgVzChHA78qEIItC+EQcP2kc
bW08HbEf0TnxvtOPwmdZnWb3Z8pToFYqOQ9NI2yrDU/MydXja0jfq1zRAIkmFY3TI+hm4ppHGvUf
bGmMaXgI4lFJc8Q58bAkuDxP7BZ8uGJd7o7kFeBG881fQna/zjhsPf9QmoE73GgFsXF3XGM6WaTX
Oi3q8OLTGCVAzZPKmiJSercuTkIIWQspbTYlFh0lEe/VSD6CFo8pC2yk2MnaGIjRjFAOxheLlpn/
Q36w6ygQuHgFCNzqzNwz6AikKqqk1eVnOkVWb6zfPijNFtZZQtRDBsGtxxZHSlC0T9vTMTm7fBuI
K6T4G+ylcAQn/XjcVnyFB6GpHR00wA0pWdp6rHFG5kcGjUPRZUdbsjDiiDaevpT8MUNRezM5Ak0f
Y+EDzjxMYQK7tn0LJ3gFz8rhjfTbC+yFKKS9oSFkLSbu6v9s4Wm5TKt+fdh2/SGFS/rQgTDxWwoD
6HognAN4J48fA5cPWMZ9r9jqDAZeLoOccIKh7G1xxk/jigT+NRhaR4vdoi3yr9eYh0ZUkzjaqfZJ
ubUa7nxutsm3KLjB9lNMJhdworwUQBDmwhPW3L9RQOl/Vjm/h7G+zBXtlErZxIQ+6yvjOTb/m6tb
kN92GeJwlWuagPvWbrLtz0ymojPqk5NbRl3LPA/JgIxTMUogGMKfy1Mox3YUWw/vTSLFr1wLTId9
TGjES+DTYV6xHppFJbg7JkvTIrE4/ElWm7yJgBY1WD7YxCDmuOwvtddr6325ToF7wSrJF6er1Zzn
iJgVQKkSSICQjAlW/2M2+a1GgyQodx6WhDy/U8UPnggslUzB5tNMvprN5ZTCqrSjVAWzC9M5j6b0
p7YOEbVTux9hdvrX+1K1P4KyIs5kmavWjHkTghMN0qcbCGSfo4dlY872GZFSyaRujJfQWC6fkkuy
vJMUSLuiYg8VSaY9Utu1bSs13GUuyQBaGLofvM+7yIoZR9UZtJf/LNGhB/VAHMT/uOaT9gfiddKB
z0ByRapov48ZN05UDUPH7Jbppe1XqDKgppLwSBC/Trqvbfoeiz2tb/gIHhSXbUbhrUdw9LfN0cMK
7KHCYXYHMs/TkZep+Khd63HUaAbAqfoJPbogprBhaBHZSmupHSZSQnA1iMrSfV6Ii0whSy2QoEN+
/g1jlx4/8S2iRP9V5zoniSD9d6uX+60L7dfcSnjSBeF/RYt4HFFnDkVs/jC1B960tsbXRi0xDY7u
CKSV/VoWJYWTLyU2oEKim+ZC87GOBk5GRIeOPnho2riTur5kI4IbmXsOQxraSLgsG5AFZ1w2AQtS
En4Pzr+7stM18zYHbsXfa5I9CFjeBbocsZGSy9nG6mieTvMN+4CnyS7QF0rmoSlolievub6vnHhQ
WhifHhUDsBNtE4ZQbYyMz28gnrvXJpx2CGqjjesN17lnyDjx88Fl3Rkde5VrWqxtk4msZkFSjlpF
EEHbQBDfz66taE34xeHxihgYhORnNN9Q3a9228EpvAN9wzxm150iyO8WZwFtUZVmkv/H+kxl3WFl
F2/AmERMcv3tvuLYcbTeSojIs9Ja/NRGw/6Em03wyl0L6fJi6OtrBqg0dKb6j8/GsRl1yia6+ZI6
qe3pSkqnCxJXV43RXKH/Kvq+i0ZBNgWobtUSyQn7TrhqKibNxFnHp+Gz1szknaBKIOoYb9/Yq5lt
GUNAK1JzaBDD5MweZhqCcoX+Arbs3rci6EqYx9hyMCb6RRylNihqVMAzsoDRaxZ8DTPz+eCaJhgR
ERWMDjJp9an7lbpYmk3x3xZFtnKkQy8L6n4TLPX7JIBXg5q+j10oji5flZWe5z0ZMVtzF/g/hNyw
hoObU+YDm29lUCN+byL1RORe8OIMvDqGHfv5Gk4Znx7wxY2c3Hgsu7HIAhSfs/i2vcms/DUiKr0Y
/AS0qLTJQs/KjA8MCaJpgAji3wMTj7bUPY6+1U57LtD/ir74qRyqdS+eOEtU0LPgP8kf7OY3yiZv
fWhZFt/eWHThpfWxJIO5fIUdDwwkCpQOHE6HfAv4Bhrb+0EWOHYQ6N/FHWEvLMsnr2XXGbRtmOhd
Msy5/8qPa4l2O+LLhinl4OoDFbQIm+SgHnivFJqNC2AnyZexdqBohlTMGwRITMPJUeoct/tpXz1u
EkF/iPqNJDCMDbpw/DYoZzJI5wOXvjGraxweLZ32vNEv+VYFr8HH9dSXgp3g4hiQyAR0blyasyAt
uJJvKvxumQm9hlr3vGM3v/3O7NqBfYxwYGi3K9hkFB6Rng4yxhOJWFPKC3HoHx64EWGaOphW7oqs
xYfEXv4dD9qBeB5ymEzUb3v31z7+Fbga3f7LQbUchpRZxueomAQa+TUKF3cEsaWiWlGdeh274j86
Tu2Gt8WD2sIJg2Qkb4YlI36B8nbCl+MF34Tdt8tFQqHVitrc+PP1YI+8ndXF78d77csSDmPFJI79
AervxvtfA4N2yNaAg5VMH1xkeBygWaGdZih/f918z0SS2XKEg8oNCr/7dQ5xB4HDVm9fYRTsh2V9
15m74K9b/0DWpAHR4ns+gaQwO1jGD7BNl9LqdZGFTLBL51AHY7ryduPIdYntz9zTLDTYipQ7iapX
pgvjPvv/UJbM0/H0BHrQ/mRZ8ZQA88pa90macFOn886VQa9xmks835vV19MpkvK7HxuJ4IVcpPH0
3ktfbhypRU6Xs/SLMPqtNfANI/1+OYuZz7z69vpQ291+pQo8ckCdKGLJN2/NcgBe8unzlE3ar0R3
M5Mi1U4PvA+VOG/nS9gO6kX9pp/hEbIhSt6SCIML/fln/8AI8cXEVKGOcZYpUXUwm4ltG+bS3nnL
WE22iXOZPtdKLKFAWJtsvO8m4B4tdcU+TA80CfCGkNKd4pzW82zpuuVZTyNwxLnmx9d20JmmuHaS
zm+0KpVSwlDl4SG89mOQ/F5Q41AbMUMH5J34wpacm4Aj8mUVe2L9STxmaanPBSB0CaD+jCKHOFb5
LtU4MVFL3hV9uiWQreTloHjnKzPfByfGoRa/Rjc4uUlPj4s1y/F5E8rXlFuAAW4u7qN8ci9jWrRi
LEuWdjpbZLxhBP41egIJlSFC8AHwz3Fwa+qAG4twzwjPqggnIL2sBSRzSAvGJ+9ye+m2dAl9AT3U
Byie+GCAHNrsDXLz690xgyMp1XojqnEuvauPogtxexiCWa8QGzs/djHAvG57/sZqXc3PNVuyC31s
FC04b5qGl/3PA19tjkdQ518wR/EIaAQvVy9Y+aZAzecTIJq8eDLF7p5tj0oBq3U001bI3MizyWJJ
zLhadH2Ic0j7xanUdkBbvioR39cRvJtKFKZT8DpFnnaGMxw/mhGZWdcMpVxVOxAVg+uIYAEo8TgJ
LPKldE2GQUkRjcUYGq++HhhmvGxMeSk9hexvxmSi47JEl3+7hlRjVeCzAiBPWQUVu0h+6x2LF4lU
Z6kSSHdIncFO+N8zjCYv9HG48WTLCSEXMcusuWCXPz976ui0YePs7q146cwUSLsf4/mVrcqVZN38
VaLe/+wJu3NnEilh1akttqJ0gR07l6pWya30SCwAYtjKlpLUP5/oF47STHVaHKMTGvoAfttKtxuS
RE7li+sAed3m2iTyP7AEoFtEj9UVPwwTuGZV/taKqcJgyZyqmAeFQYENIKXgbRYW35hIxyL0PjPz
4kHeip6Y2HPAFJDa9akfbQFENXSXjs6/V1BXVMT+gMgu8y8p+QY0hhwPcHbBmlE5ejGkimoeougO
ANOu+zaWLrAyQ69C+4N5n57cbP/9hF3sMO/qLzMlOvOZKDO0/lhMzg9uanAsEmahC/5o9uws19UT
9Tdlm+CqJildE6MyWTSwrgoiTk5BD33UiIexMf5OIRgSyJmg3XPbWjJTvZ78FVNqCbS/TZVNobQx
z2j5YpqesTKqYLzWMhIns8S4hYQGGJFMlWvUCWxYPLK5Q7hipx1d+HP2LHgjZnaCLntImEfDSzMc
B8jHgLzw6fRLqV5mOJQPgw5/ChBHArAvuz2DCXdtwpbTv4rOleIEE3IesaZ5KwpA2qhNZJ3otgWF
VYwkXoT1+Fxc7t+4XSLBcyjeK6GNQ5SuoQw1dOKlFQ0kdLrAUXvYiugJ13PO0RBtho5pBio9HSqA
XmVF7a0BiMGhGVkcbcj2NHEHydIFCpevtKbrYE1yveQTQ58ifCsBS1j7/VG3LUj9Ymv8XWHBIz4a
28/D3McJ7XKRI2BMrmW29yJ5tbm2wJZa2wTpQEJrBb888nGMd01IV70p+M9IW/aAeNgWXcMWP5yz
hOU5CMMONW6TJ0nqJWDbMgGE3s4ZCsX8/iVz4sYn4uGBvufHQjR67CmGahSzcokb5xSYPpdMs7Fq
izaMx9eZhLF/0mAPgmX630+ZTgWjC3iVtWi0vkJIXVgAor+k6hP6OAgRk9VvzXRfYRsBs4Jhp3H4
6sfT9mrdZ16N0OCwrX12YjuTlaBvbL9FYmAkaXDuQn53fDguK9ST1zJ5/BG1KXkrs6DOaK6Xombu
ytPjBC+QSIPcOY6hTiUZZQWpNVlRW4Onxlv50b3r5wqfHLEx+YG5hGYNjSSDgmx5MlkQ6FmnXyfB
F+aVaY/vRfatS6NQheZLEQmP1EdrJ/ecvckNWBFnauq/4HC3rzmMbhdSEpt0GCaU6SHBm7tEy8Va
TwkznzCzCOX+mc+CGf2C3wVZvLVYKCoD3F4GngES6fgPcBJ5u4Y9BMHDVg2UVlmlEdLArW7XhfP9
WzPD0MybYsWJfLQebJIoIwp+pociR5FTQdKomq38eoo3+ad6gb6zK3m++s148+2qyXX8qjaPzLLB
yK9vc7hLIMTfVviUWf6JLqXYdJXGKpnQMC2bHBMdAZs9MuU+vzQv2FgLgG/ECkDGucMF28Nf/FIv
+Y07zP10J42u8DrAceVL7ki9l9uVk/PmkfJYGgwBtCW0ys2fNM/BtVummK5LyOoWtyMcJpi+hwH5
gOJKu1DleMZh86MyEh+6Y2R8xdCqvHJ4iz/iFlPCSrxHy8UtgKi3DNemqbzva67xmG51Tl4kRsgn
vnnbfKwqx10kDOG5fx7zftu9ecniXKkmghmv52J0rb7A5nrYHlmQOts9S1RPlsbjnXerEL7Y+MWt
Ia3t0GNxPCv2cwSBO7ty7v8ZlQYeVBMteGtsgGxLOtM8NjCPZY4vGIL6z3gpm4K/SuamWJxd9cO0
s+evVXX1s2FynkWogYLhpnP9OhC/mf41h1iToA5kHcfhCAnPjyhR5iy4dkq+B7crvr247O7yymZA
vrUjMRJ1AQ/047V3/w3Rl448ccEMyDrDQjOi5dtrOPLcWDJEXEHLxyqLPE+/bT9ymZ/vHjxzAQpJ
82Rua8gO2n1jpBjjVcxUzUUr8hKYfGTZ609qvpwMX8EXV2sSfZnxg+vfa+B0lbiXdsLRustltQGD
AO9LNzDkbW8sIN0hmvspFW5zuyAFWa7u7+R5QLKVFTvdD32QOyNx0N/Y+pAyX49trsXfX95AOgst
fLxOyQcDTlA1onL9/v6MIwDB6A5SiIw0ofmp6GV4P+X3eZ/KLzqemRWva2C+ZABoRA7a3dP1SuzQ
UDWEp5iMs3Y4nUFdbTsG0jn9+FrsFRIHuqMidp/9JsG8dO31Kka0dwRoR7kqu9xgac2IwArRgHma
eZUOCkbOrd8csuAyLXfoMPL6QRhVkmnnOOZd6qoTICraTR0n+u3fEonK6cP4Ybk748b78vtFwRMF
UQoetjU/P1fpEnqJDg5oJtaMJU/Zc/XFoQCXBh1bOaGdWE0W1sPYSe+n8poGpJKpZUuvC4l1v+Zg
Sb4EHvmcZP7C5lX/lfQihVGOJWHgKzASW84T9NYeY7jqQzIezz3dzPIYP5Rbt/42mUYX5zdN1Qua
mQPO3FRzkARqvYRP1OiP4MU8jG2PaGVugPcOni3xFMyvFw7eqKsJ5HRi73smdoPkFkRa0TH0cNud
w7GSQi9+UmPPXSIqU0yDjw8lQJRNJIyBbmak3sWHpEC/neL6HBUwbYGGtykMvO5SVplDQPUYIjDx
ZIbEWE27EU0FO5GnlpgsGvtpZDt8IRIbQNPhsNaoS+qFBnrxySh13aqgjMmi245I4rHATmnJ7MAq
kWIH5aGCTPrP5IwNYOmTB+K5n2/1yep2CyXmDifCGQwPXYmlRQEm17KRl+SlslbPegkx/OLZONgF
hd8LyP6bBrK2fSNgzn6qhy3UWkC3xYFnLdzJGrSJt8B/v/n27fn1COjC2wh0GKof0ha7tsbSGmwX
z9QfeuEpo4LIjrAg/YCRKkBw9FbEFSbi1/t7FjLwmW7jtcwnOIbm3xBMu7xwMRn1+yKSZ2NCAGDk
MVsoi7SG/Xzvh/GE6GJqULag1sB5C/ANSVJtG2MP5KTgbAfw0ztsZKZT0E+aLNpqZEr7ZIXNJZZW
JtLb6CRfmJLyGz6hjYpQg3ymjr4JG+C4rVQ+vBbfzoiVI4SO7EY8SPHD9dhMgvoBJ3olhL+i8fpE
t8d1KWIias9ZutFvWCf/4CPlipBboBsjiEvhmaCetS3EmC7xgg0ExOiy+Ya5BBSDOAPldaA/DDG+
eRymQdt7H6jqpJ2+NtwhnP4bH3fHEvQBeg5sqiMTdQipZjzQBgulv1/Fs+O/Vao2aHhe1rt/r2yE
Qvom7vH7aLK3iEvlOSfB5AzRvRZb+WJr6kUctBZHPQ012OIxD8dq0HzHmtZfIUgO5+GXZCPi+ab2
1CxPVr5gnV657WSRGx+On+LSGJJIIHHvICE2TXX7B+v2CBKul57Si9lsBB0BGBVKRrgd/iyoobSk
AvvvSj+m/NJ8rlJW40mjgxwuGaK9nzGhta7DK58xS3+ilfIyvMcwR/wUBB00EQe6XIxYe0Ql1XHD
aIoL4V9SRJTxmKnMTyU6jaMQGB5OAkio6hneXajuW7+4Au2x5iMRr5gLejlTm0ctF9ODFKTKj07U
zdmJVUNAlgk+lWUXl0CNngOQRckeat1GzAlSock2a2/qQbxacPDlqB1c5aiRU2V4zzQ51lXgRThC
XoEcxPgCTQS1P/laEjvl1CUktbiVVWL4wm45WU+pFyvyu/pdKa53KxgNTgjYermbjzW65RIHhrX3
/9sbmnqtCU/macO855yw0WlnuQWhOspRyw3yiClJaBxI7BmPmp6pLKIrjJzGT1jdhEK0pS11uYat
kg/CtUSapdw6Rr7sxIgQVZWthF1wbnnRSuhEUnIDqZo5gURbyLMuhviDft6REuKEV2y6BRLWNteD
fVN5SqFF+o+3yVl7eohoDpXwFox3ifelF9nWGXH3TjsV392dCXca3FEA9qGXA0dBNjwWuVxxpqLd
a+xAuSqEAjy0BJb3kMuE2VrVcJA1gQA9PtH9BKWuUtc2E/+cC/SUYZ2KhV9QFPkSPScSY6e9OnU/
+/Q42cirO3NtegVsi10BTH9xTaslAYbPlgJnw4ICO5qI22s+hdO2baEdywCDln8uB5KVVknVri9J
RvrUAtVzYrw8rztKiPs7gl+N7AFBIEX8jQI+NTpRlzbpeYDfZDQ/PzK4KOQXpYtWen1mbu0acYVD
9B9WJT6GKmbKh/jHC/ZYXw3ajoIh3g1gy1aKv2oUW3gFUmLGebBveSOMFFTvq+5MfIgRf/KN03Jf
XLDqbzRNcifIhoKKVJpuhWj6nZoh9A1wUD4nStoEXvYrWEzZR58PgZCJB5dMNSK6aRkDOhmA5lmF
p7keqUWCsW+7q/39aaZAXJ0MIvng4y3ZMcRRSMcWkjSsuM3vzCaaIqYWqntafrI19OLBI9qE1qiB
zadUMkQjWaHXejod2iiivRYOXCwrGqvaC2V9mdMRgtTO4ZOIjpR0d8Hi29/dzHesbJcxW2TRQ8sP
1wUkGiHdlCx7353QLaPKqprFOWxX0l6KyBOLKREQ4QLUVfQb5fpGQ8UNKqtJ1E6HcBT/ih3+dTww
NTkCUUrY1Wmqe+oge8YsIBTr6cyVXLsNSDc/SI35gb9KtllcCo2O0/JSxT8PJa2f5RT+iEUoR+2u
fWMEaWZtQ2YmpCD5xiJI0muaEtCRoCJx2JQpsONWk8cxlUyybRc1N8jihphGl3h8HHZd35020rG7
1zjt908pfAuBxB5Ic51oZ9MslhX/WLCXeQROeF1JZeW5DNPySLpQ43JKR2/8j5+4SJn/HQazEkHe
BQWbnUcq8TWFRflHnqrQcTUAZ6HTvXKB/wc0oZEXK6bJnYjRypup5RvStv4+ZU9sdw4nRW+7XOZ6
xaLY6jCS9eBzgLurgeS1KkDslHNN2gnAPtAEqC+iHm7tdW5LWKzjD16/xAB7GrB981+Ypc30bFgR
4IyWDsSU+aqlhdwtjolJJJ3xMthTZpDLqZr9Cigv55b+6awC8Elvb6FLEJIDb6+BYSfi8kM1Jl92
uYrXY/+fAisHq0AomvkFAMMhv3lXBM9cqPvS60mxiU79kow84woc/DbY3pI5cim1YINDMuQf6Mou
5nBssB8100jYS2fs0Th5sDal4q6aslf4fNhHjyfEBA5sutc64KSK4krSyw8CgbeWW3oNCn2yvIxl
4vEyL4tMLyz+1gdYTiVuG3+bL1yH6jd0OS5WIwrAHLXpovyFZrQfVOH/EOQkqYxtABr2YmGz6+Dz
XivuhuqN5ytvNQGp+8H/ISwLRA15gvfe9wwqUM5bsXf64vljOQ/cUSxz/boXvJtu4A07AgLUiMuf
AbSVNMososR9aZLlb7dlEoaSCroyZy0ac+i6hGxXwo2Nk5k852g4HmhlQaIQvLC4MqgfmC5Hu7Bx
ik5fE4MjP32T5vhBvRsHgtyaJwVWJ2NxL3hpWw1GT+WcyzGPf3ZnunQDge31Z+jUf0+8ZcoM3w6s
JQFPC+11rIMwzNeylhiPwDah9JpRiS+wPrvugf7np0Y/yDItPzPJ3lhrwNWnhKzDVYRpOZMSDnZh
64/xS4y5vr0ygLEfv75YSbbhLYjrakOSP2Wcs9trI7yhKA+4uMyGC8oaR+6wBDngcYEgGZHzaZu5
6YOzH0Z3BWpZ1s0alOr/QTwLgQvSVNJpTsWAj+lNbDmfRxiBWXRhnKeSYd7sZplHNVpgC59+pf6F
5SwIKWFo6SjEA5mzVfbnMWXHQfFda5bXUxOtYfKWZxuNFknWxsq9qyl+8Nl1/9vQijveCP9g3V3y
sjGnaEOnDtLECgbATpUxgt6QMauvNqfKfMsItLemM1Zp5PGAmEssIEj5brvi4XEk2aAZeTevPJng
GI6hPXc9ZJWIyvyaFyQzsczF32wcVICU4Ng3t8GuRtdDVUOfp7r/lmQODl+sefVgd7JcXXp2E0+b
msKYd7cMh1QjbYXaY6QbcPY/gS99rvJVmNCecMAjWfIFWfSPKd5xYGQPyZY5oSyo/3uHondkW26R
G1QK/8b8KQLV5H7leFdtncqWdCIEl1/E+fIpMeMghu27GSGNcmad9sN/DFFdrfRNUjbKOwrlmMW9
l04ah44dWPobO6XBmZ2+YhUhmO1GSBZYjxXKYaaI7ExHs7scR6tr04uhxBtonuG4osz97tJ89Y0+
OQHl0CWS53f1lCU6l+l2ihOUoQZ7IGmQYsjyIsFxR23ym4BMaz1A8gsyiS/aYYDGtPAlqX9tqikT
yWMGOKl2stuPWavs0xWukUnID/veVrLC1+3ZPttBJkN/yxJz0LLoQHpQ42rMANuLQ8SS2k0ckkdZ
HIlodJql2KuQQK0AgyZeIWytYJeT62QDNj7sWtg3HegBpkhyQZ6B0aW8ZG9NF8HQZXWHwVxXo7ww
ZPBtZUPtvp2KOzVBULJa4+Hj67L4mJsCcLdqFevR5WMDd3IAMy9n+Si2v/h+a2JLEabVvh2xn/Lw
egAYRHuE3bYX9UFQmj+/mzzWpmObwTvOyuPF5lqhNz71oIlGY8zKIshl8btTzx6SR/UQzjDxvT8B
nANjrDI1X02OJde2XxOm0wX+9Gw3h5QSaJBq5gXCzcPHMEwUfU2nBp5WtqFEVP4RVRWBQww1ND5v
RtASvLpb1C3w+HUTmur+TX7k3Vons+QKG+XNW9hTLVr8b5e0bQ7cfH4j/3K1cR1OlKIWA78tXoN7
PvOl6nISZ1NHemnZszSokY+7I6pznQA0h4yf5iGF1rhW5e3oV2YE7zapfk56ovaDxbWsXWM2Y2zE
sFLvbSh4D9Q/v8+bhoFatvD99wxGHx5sgjb4l6e7aZEM5ddhm4WF+rt1mdbhPVtNSX2gBsvk7ngZ
JZVSXUO5LgAI0q87ghuPDFBLXKsfOEFKhFKRoxy1GV5yT/YDElHD4DJOcqaz2aon00JKPrdAIZ0A
zO4klPl+20Dh0EqR0xgBcQQ/K11eZaD3vaxHGPoPTdT4Ie2Qf89FjRBeRse0PewiwH6b/HkZNUkr
I/xbm8k3TF5BxeWcuG/Vtf0G9cI3a9IbEy2qiudYLv3HTnROeQElVzUNbK7UuzF4R+enzfqEA3Xk
nTxuDs3/+4HbYsf/duRwiBrmKs5LDRXOBapRLiR4S0KuGU8IXGqK4ATY7ZRPjU9UBOp8cRKphGEZ
ukrJspjNg8DIHR91aSau2ZLQFseNiaKLPiigHd7Z+gFVp3VayOSgl6MfwPOZ029I+GqcIpr151om
qWpXDQIGLnX6QNXZsmDw7c4wpzXZRMsj6zkDdrLyxriOMgs0wml5etu2x8A5NYKZAUQ3/f9tFnpV
ToD1o5fl4dreR1VXyfGWJOD3Dua7EHZG3FUD+SG52+WkZNXhkFFlZxzkK970IXhJec2GPOmF5OSB
xMT7OOr+f1PVVkh+EIekZTAtIPnYbMbKkZysdItbbGFhqa9Hk7zapiiRoAKDKr86bGkY2UDpG6Y4
DmXnM0eAJD84XE8mDcHxSo4prES+FStvJ84AJ4fKRZZl1GJ9XBLaMpUfhgRvQTNTd3ESxG7lqYNq
YuFu8xL3L+g8kODORP+2uD4kw17SdshnwhijNk6e3scVqcYc8qmNFB3Hm2MKTlWUDhIOBc6T9gbf
mCnlwUEWianEh6HwrOAeyyFyZ/IXCU+R2hHDTJVQLtxTHOaEVdJXDPOLocbUl6sr+7LSJw5K9yTL
Od82SWjlPGNAGt5wWplGlbUepS67LiRWorou9B546ZYp//9HHWGphNWiqHKqweJ+euexv/rZ3XZ5
IbdoC2UEgL37zhQcZMzL/Tey3fRFvbhgFHpnkocvU5sZa4zAC2LYxbzh0S88NwSHvKLfrxPDVcWp
dOyJk6PEg8hAhVNFPkJCNrd5wSDbBrfS6W+85j0Sd8GfEt93E2EriaHB2azcNp3anXWvukGMIrV5
6eYZA2TptCefcAGwVMfcPWLexxK/2uskkJDeEevZRNWH5Epqh6bebCJL80bHsRfobx9nO90gwfgs
6h5Vesf/mgJP6cS6Xrew52z9cbnn1VZ8mSRpoqWpSumrIDeqqJ77PEocBeIrcq0yS3CqlvLXT4pj
FIGKXpBchQr5AP9rpQp6LYtRT6mnyw9aPxsuQx24YuIAwN83oiD2EIjfw0C6Dh36LhljG5KzD8AU
y2d3UafKHg5FJQ2nKa55MnRcRanWJ9tCxYPwLWZCEGHcwu1auPDGvZpRE+fcwcDExNZjyuwDKjwZ
gSBte0n74DVH/Lqvc01WbPi0wtzlJV3Mstd8Pvol3r0DiwOKx6o5tC8zYDctGWkVbIuKk7fxhuic
6mFXoIzUwPhvwXcykC8gvdv+p9K92xMjiDelvs0WKjntrm/gK7WQ5GXCdZlWCJMxdvPhz8Ys2+XW
zbZ5iMzQAbE8UP6GhDxoK1DhYB6iZ6X+l+vq8Afg8tG6Y2AWRQyCERoH7qCnCvCeX1TM8igG+sdQ
XrFwv2h2IRguo30eeRMRLTyFOWzA4SNuKvx5fjftAFf1iJRfW+DqrqyiA580JCemdmyJfsBs4nss
MjEp0O9Vj0WusDbmOa/rvqNBw/e65EgS+H7eTZIwzY54uFy66cIzyrJKQNG8l0zDi9CeeWffZuHj
rYwQnKOEd/Mb/jwuQH/pyrWrYBFaUhIglRtVlCWKt2GCEqGw9TGmIChyovIWm7tspbH/KaqNg7sp
3/iq1Ccofk672+IxIYWHtL4Mamt2b3h4QUIsDOxOrxPpm07JXVOIMfeXjvfmayZRzepqkKEUEG+5
WLQX9YSkclnZCI187HmQjqRZtGTXhDSyWwUhKN0yhwy6WHt8YvJJlGOov4iwyuBJh65lhNbOae9F
/pH34Wu3RIhJlggofjeq1rU428UiD4OV7jDUfT+kRodb2TMhv2GO9GzvYIIswXNsrcFMrdFnW4N3
vahMEriU+dAD1/8RuOaZ8bdnVB5kW5dc9LfnsLTjZKp5m2aIhRqbgnwr7kUqjvCoPvr2hyVjHWQn
tAVMwd9pmVzHNcy1IqU67h/zCDWn/7Zal5966vYv/kcuAXIVBGtRcH+Sq9Aw/8VhMLRwN+tqfWgG
EszvwWcqOVJnXz/8qrqDLb8VvrV1VPcFZs11PNHdbyupUsAo/hhen19dDjN+gY3S4pjSQJXoomjV
u7k2JzTIQCmZQM+C3s37O6d+MdYk9Kv4Hl14rEk9Px/45SNhQFe7pbrqtqveUMjIVrjps+oLt63m
zzE7JHSpbgdCmITeucbsYM/OIUCiXdszE43aUwCQteSYuS7jqBmdXh4MVaNYburEY63CM9kim/RK
swXyfeAlc8TST/5RsQzVs7l8Gk1fJq7f8LUAJPeWtsQZzuVTDrU5PtnHf3Jon3ZTNdBq0D8K+idD
ckXkv4T09OBtb7nEvqjpt7Iqq+5AOqcfesuexmg9ZLo8QLFukVgB/7H8SLp9TTdOiwIGhNy3HV5O
brixRDmSn2dcksMjXs7R092vNKYo5j7ue/x+JWfANLTJDCU6ca9taJIaboIf0kIE27YMJTRp1SB0
qZ3tfm1n8ocVO5tesK0nyR1l9+VDlfQz19pxIuE4yUFzqP5+E+S6qljAf7Z4sNidSc/wx41Tzw7R
WlhcaO8SREUzW6N2GR41GrokeNb9UtdM3t/b1lDnWyrwC7DlEMaSHXVkKsJhjOBmAypNgbu5nCPT
oKLTAqsm7r4tkY81qsH5xuOKeKLBHB/I5cTCTvtISvhs6eXT+3+mNP+F/PXPFGYeRF4GYJd3nOV7
gGo95BMs53w8rjGIdIirrstYiId3/8Zr9kDqXqxnLb3FAASJEuonE4zwIBIkB8x2EYSQtVhqt4xF
XcBLDdd47/d8w0h9Rhd3UQOxKxCM/E95RL1qb6v3D3hRpF8wuky05WjrSwJhUlu/+etbN2qXRRLp
dYaDcIhDgMp+s0CPdq3bd0Mu4KQzdcw+ZgXSvDOu/UK3634qkdJGshDqBOKxQK6ri45Ac770GAA/
1zet/a2wtn34Bwa/i04giDf9fkryOnEDqDamDcqBLQAdCtwWPCxgFDoUh2yb1/ZpYwbrbQ6MxHsG
oijPrZwcE4TQviqf5B6F4GWVDBrweFCkPyJy63/wzno9qo2bbDXXpg6+QXPNDycQQ+tZ3wUSO2ZA
BU9o2e8BbWnvSQcz3a893mjqNE99w2HBgR4QFw4c2mUzWb2WgcyblvO8smQfp70i/dAnSe0y8hR4
HFV1UQswSrqIsejyZIDZIT5mLr3E5U05HdXi38MafK0f5p73TK3ZhuOh29UGS1FOjZ8WkzBAgnJT
9b4RIJNWsSC6uJCtOeZaGbEcr55UKrwrlSQEWklnK6c4hCA7P43Jiyfa+Zg0UIs0qQKIlV1GF0iG
VhNcX7008PYg0fna8HPyWssF9XrZP6iI1noPdBY8kxdi/jR1JXmo+3cBV0eaOZld9OF0DoYFtREb
Kvvz2WCCklLMhJEmFhFsPQ9MY3NGkmEDC1QNNG2SUkjbcTCTboF6B/l9dbnIXzMDQKOUMtvMPNdl
NCXuBVxoxOOA9H1EFGNkb4Wri/fylT86Ys2q79bV4NEflKmN7XSVjTTiLjzjHL26LT9HxFiaN1mg
9sgRuvaco6gV0dKvTsMm/5UOaOTmtaZlDjyrqdPl744cu7RUUTQJEbMQLDBQeQT0cbYDiNONMK01
VV2vGCrHAzrtV00H8u1VAOdePUHAKKYCLDXNk2UwpHxQrhEhr0w9cskw1PfK2dquuSXPB7nBUKUT
u1SZzfmAbzBMmHrZFYG2xcesbOOYXQTLlnwCd9lRpNlAa3tpkLO1ktl920H/uIUnsRIhVQNBTvpd
xomjBiaqnD8leO2htQ3sOdXHgiJWQeboI2HuXP4rJ0T+k3ApzPu9VtZcJJn/nRGM0dQYemQj/dBV
Exg177UMDHEQ1UtKF72ZQV2mA+pgW5HkRnhTETzpEv/jZJ3DJpRrDMW4pzaPZr1gGcFWmiNm7RI9
aSfdQzxjJ4ZvIckewS96uudJrL5mmXz24A1ouLe8l1e1iQu/3KHgwO5/GNJR09XnUeRUjd8PRQL8
R8RtCjBiz6p4uhBIkzVLi5vZkUgjNTN2X3BUXaBQ5KHpwq6A42oZLMZqRuvrO8i9fhyO7MiROlPq
bE2fMRnRuirBAoI2m3p8acnQZ3gPq1HFvqmRo6QMvR0a3IizgGRMNOLOSnfdAg88Sm+9vLnVHeye
JM4nfy6A/Tb+mDI+gbae6RBnVEGNVA98FpPP8XejldFMc+XdoJpcZTRKb7S5s3UzaShf7XS45p7x
/p+3kH431AjeTWGm+WY69Zs0asoLLBIpwFfTa52c0ED5Ng9y00bVfEAZE0w2PghL0C47ixOIYIsw
Bqd9L+IBkL0arS+Y/G8AjbZqMxySxbSLX9XUY5jaT5x+zFzsL1UVXqo9jErapb/UyTGjS2otRXjM
/amxt22SDXD+wfXQtbLtTYhiWP6T4NodaEcf0D7oyUgCzXMZjTOhbDJqO6IDh///WkpSL70n7D2n
NR9bw9ByLNj6sN78jwyBuLooR6DK6M2ercB5pI7vYVxsDc5ApBujMONazx9HTWUzDcW1ELQbx3DG
yOOrUBZW5NgauuWLKqV1g66oBtu+EtWTljuTzGWOqhoc1XRO3VMBiPyqQ+tfWuIdPUHPNezg6uqZ
4ONFHRF+KBxE7dRnJTLDsy8EC5tPKmwc7DrGBPjtMNpGZbywK8WU0NIjes1zmeqa0BFaMWNFKpaK
4QhPikZgG3EGShrsu/dC+BPqVGKi3M6kvzUlEOjw47SQ/BRml3u35o7r6KeIufyUrEoP7H/wQAA2
WhshsLDaWFK4l6QJzO77O0zQE1rMpm1ZRYLZT426SAi5S94N3cfsYiKdzRFEN6maIHIfzV/hROX7
utaFSxrvEZChiXwOdeqqk3r/ux2PHGaougadbrOT6yBqL/pPhohyTRm9PSWxBYZLSz6oCiuzTxWY
AU8D/PyBXmImfJbAOm7JhWerHfAvwe4fNbZ16oii7MrWwa8wspjuXReoBYP5YW/yP0OAk6EQpZVD
pqR120qFt0FMQHNDkiouQPtJS9Ojxd/TFPn+VgrV+MwXEtRyxgInJZCI2bZfTYfiyDMVI4vCvRCT
zLl1gJvKlHfxHl9BQVVjYQ4rsv4kjX+N4uky2x1Sm/F5GJlHA0HV0lo7+bEfx+MnQgZkPo5qbkSh
gRw0fNmchO1uUBAXy9P66t+0ZFOrLj+v45TOSzBbiPjjrXfFUhwWnSHgBG+MWzxjtst7XlDXVlK2
jAshIjCBpkyBWCigPTPbtMKPnT135izy1XMldVBvoSQ+JZdaR3G51czlJ+iimFF/UIPrK9zBNKot
E8M1K4pv1S6sC/9WPsozJ/m4qK8o4XPfBIXIP3C3RucSWYtnLb2jyd4friARBzQ0yG3CNiT2o1+W
vrezFIfOhPp1DxrDdZBcSQHy0yp7wycYZYpEbnS+8H7mYDo4cNC7UBCeOvl0OHR7hA1sm9bXN6RQ
9DT3BuBtrnyNIOTHS8EyiDiNW2k43ooZg64Mku/N3O7JugnoHXv5UBS90aoXKelIRwXJBCVBgpUs
pzg06sWGHWbvompdi+DERyfb3Db2lZaX3SmjO2igOsuq/ffqMzA8YF7DK+YRpZpoa1RB7gb8TL+Y
0cj8avdnjKukNv0vLIv5ShCy25GCxEwWvZVfbB1fmZRa1Mnm/pi+f2qWgVEpG5zfLL6qz/OZoZ1u
beb3gmD/rcBG8BplcbdhPVGGH0gwvMzdYJqrySNN+4epS0FHHJeVuOOA+Cr9ctBbZ8qxh4Yh6/ys
SuW0hLG/U+FxOyuAjD9Tq2ngJecygVXyJJZuuX3SPXGBirpIuGRXeU7S8cFuSjFYvDVG/aAiRZzx
kpL9qD69T54R0uqok5e+bY8Mf4rtt95Xhr9J4paKMRENs1Q634s5BQB2TNFEb7z2qtnjL1tpOKIS
SMx7Az/hAzZesr3YAh8z6cAHv44LmKONNsM9BvznRdfc3Ww02duugoREmDgSzqGr4FJXEIKh1qrf
NklqVeCzX4MIBWWJKakkv3FkXZ9s3HT8JJIaSDaIytF0NPTElG+CC6Zs2hjekGqgg5IHV9B/POPl
QE5HV7FTgSkemHGa9PtQvD3EoR0HVPrnVNEz2LgYVvwYEuspPyMTNqOR/G9T5SIuVRS4C+dF7T70
+7Q0bcF2YP8JEID7zSRPexUR1qwgHTHDAdmtzi/m38D/MsJBe5BqhsHct4puHfCB1KfFExDWLRgT
CDp/zRtc0RQOBgWfvqGHKA97UzYqxAn8Ig+OA2cKT405q4ZeqWOFFHE+DN7AjJWtYNrz2wim/+xM
ujP7qbSML5a+kMm9ZVdks+P8WJo8zaU0Mtv05Qs5nYY27M5c0Edj42KOoLIyEE7V46iIk8ueasRO
8hEB3a3fenxL68QRfW1ucBDIZbFjmLVmM0D3XGMpMmO1EXUvoWOshjhKLbOnUYDkMGMXWXfPUrsk
5h90BvmA2J/dL4GWfq2L2t/6Ign++rlMzZiE6n8tpdurWMs5281tPWzBZEJnLVc8ZwpaDi8ejwCF
zqpPLuRM89bB63k60j/BJxGX0ktrB8OhHSGhhY3dwBSOscKLZWi0F7aB2+wiTg8TcJZNDRFM5p4a
DIxpKquqL49OGQLg1QPFVoLVkQbRiRNwnXyVNv2DYMkBCh2sbeas8EV9ZmlfEIzvmBZaejjMNkUd
b4ZEjNWK6JkjxwYQyJBqMS2EAQ1DWSm1pj/SnJjiDhi/gFeCoZD+2KpHPy7tky9Y2uJgomjtqlZz
znyS2tJLQNCNPEE4rHlFoKLb853xv/is2BC1uCB6a4UShG0Y6hqDmNvJDTEWW9gY0z5WECjZBzB+
znSgLllsdvUOQTYXp+zlBIbsfdfehj7r/+OQnvJiZEIBI2AUNILfzGv3HqDZ+it5pAf6rrJ/SRPy
5blAIXzR9Rrb3L3vmIsNR9h2/eFpQMV5jXpTlzuLEs+C2xko9DB01wZgGDGptdu4NW18AXzTgtN+
F1LGEpHEw1aaJWIL7lXHN65cfTV882Y8mKEXBeqeqSuMYc2kQKrxSaBuH+jacNNeJQUBsGV+x/tu
tDST4FKQ0iQ6wukz6u6ZaZFsNbAMImSSUUB8hAko54l9aNZ+ufWFOOcF4Kizs2RuBvxRqidlxosW
I+hYEDOa4WzwV3j7RYq/6EKAyeOru/9hcgYJtgH1q79IizCRdp9M5s1wrwliAbziNsthiyKRnx/Z
9kif6rR7X3Gn8MirqUv5ZX/NUr5Zu33hUhg+lT6nW1X46WNHq0EGCQeIwRs7rWAuoEBDk4qw7oIC
W5Fie2HVcY4QfrQi63FhrtmQcMCOO5G9FiHPNyOlKHXaoBVg9+SMT0SL2dc7E9L6iSVL8C5cXv8I
BNN7wSgz8QES+Un6Oj7YYWow5tfhrNegSPYLS19RJwmy8StoA79KXP+iVJdBWuG6cKJ0n57A65Y3
5t5tBWBfD1Dkbma6wjHWnR2xx+bKbjq0b6z1XXQNRu65ea1/F1STi0B0Ur/+5MxPCFbWolw/XKjs
ifofHNJQbXs8zjsmcjuKKRMieV8T7f1Bn9I+1p0YUI1yvkBLf99hcU7unXM1AjN/GOoyBr34ZkWO
8Y6yfxqx4kqLs/WXNMF6nAjuS2JF3P7uDlWbtWOYXvuyo+gyVKhPcMd5qaVOm/1TBjAEjZG27h5k
DDNd06FJJqn+LMH0D7Shy5CHcLqfSVqOjkVyOieCCTEkEdO1iozFtXN1l5JaaKMcKVUqDKMrD+9p
oiHz9K/fMcrVMwBFChsWqqxZo4kZyL9GHEX9jbpLZLwZacAVaGLPSI44NTBLVnfztBOdDjBfrUyo
XKOr2p28dvpDXQ8JrsvA6zZSkgXglPUeKYedoqxlE5nkj21w3rsfyk1vfBBx7f4stQ5T0AMdIG+y
Lar6cKLjok7MWUw+CfqqgRXsOROF/YZZymhWgVbQFTrJsr+GfD4szHNpNsYqAKUTnheSUxBSfCfl
YrzKitp4gAzAxXLLvrDETiGxRIfwSzxjePbh3DT9X7LCgaDSOHCL+gEGgnIJIuvfY/0SoYtes9sO
d/q1lydBMan3q0vctlcH47EXSuN3H8wag58sT6ckSn+FkJXSg/46SZxsfQ1gfJlSJTZb6q9+teae
D26u4tbX0kz+XUgs0NWk3TgfiNRph/vPIvPQGHWUjZRHxLe/vDVb0eAA40PF+nvdaGVNumGlrCgE
+OLabgnrWIa2Hww4r6IAgA+uc+tUTt8XTFqivX9p4aVN6ozykQ4gO2ffmgWmGxJv/gyQ3n+aGGjm
m9NG33e7e9O3dPrOKvLoD6jZX10BB75eQtyjE6IAM2wj6U7xVMzH84afbbhqXWYpjgUjUxQsQCXN
01lQk6AefQUROZvRrdaTOnkEsivIhrsWBIPl7xCVEiKBDxFjmqvCxQvCDJey7rVVukZeAnf0RQ73
IbC5Qax/zkvlQaZmDPb1oQeOOWC7SJQp+iayqWZ/seM1DbgmgQkunlDsvDQXlrXHAPzXqqxpNJ3w
7YCs+/al3mwyMXkQPe3/6fHHJXizQNFlGYCfQfsX5rHabRmwFtbSnvfHQB7Whz6pjxj1Fz8fecS8
yX1vpnMtcGNsVkN1Iio0Gp1/idfNT9/mxw5RIIuhfZDz/WG1m5YyszsZzBSGrsXOq2pjiSf0WaLn
Bje8Z5tel/loyG3gMQr7SHshkOTd7PygrWmLxZu6uaA0HUs5AAcAvVn/GYa6it88MbaWVGcnI0Nc
lypiRiY6vYXy8uIYBtCzQMOLqlXEoqDIZNSaYNarxv92fuds6ZKzDUFcdEHTvcUMGdUN/uaEEcXX
CoIee9oGST7ofsl3t7yQaoEelCpTlVm73utOSOELeipqfK8KWwNa78u0ysJCuKeX2lp/OVgxjdah
WJMDxFl5VfqAdTM7PBceGWIL2zhmSYjRsiiZI0rpS1ne6at5W4oavxuxeyiBfWQ6cIp9I1t1GNKr
wgJFWFceVr3cGjIk1HjqWKN4TpBz0pfSW25kDqXjtmslCzNWn3of6i7TiCXeyXarsxF6h0hwhy/k
2cltjj0YZRE9uV8JhfxOc77L3vGri0RPavtDmv+lhONRI47UDqV5YKlx7AJhIMRFFAk0liZmV3Id
ld7xsO+/TOBG/4BXKrE3O+DvZgabu2r6ZY1F4AlCgvKwQM+hE5VkY22WIRSJLK5CnPrLjqV8xxDi
tFdwx6YWL+CUFdCXurQDX5ldMoc9hSCBQ1BtqzFh6rZT0MGDIP20AVb8WBjIQglWoNgE+bMANXUD
CKmXk+WK/xH3dAZC03YwFDrXQHampXbi/nrUyeR8GfCdHAgVxp8COWRgpap85yEw3A4kdl79eNH1
9YxSSVo0VnfM96/oVUVQu45xoJpkTrpJnexBFFt1BZX1cydJcvA30sYPiCwe3sPnd9sNkHPqREVf
6cPfY5HfRMD4hehyKNzNfBHAQnaButf02/kHE6XwGCvmRImmahimffDAw1w6AMh2ITKuNTQxUi20
6SNAJ3ZNgY/Ujkkr00lKQpQxjIAuAsfYqvn2ebbdir10MYqxsZrwwav90mnPGNAbKtS9hdFkr3oQ
uARKvqqR+LBTAO2GyXQ+gYzHfwtokgtCsvyqcZ8GrspgHiaRiPS75BPMaCNHA3yI2CmmHNxJUm52
Az3r/AyufTkszMLaNHF32gi2OUb6fkvBJFVQdgOwSXax2I4BjZWKdDB1Gm5ECKA3sTPDAfk6fHS/
fp/glCaTJeAkXT0tXsWH1KhYC33SnWkmHz+r/T+bOVpFC1NKqD0VBZX/2kKkCCcOoPeZQzqvzCiD
kJnNgKh9etCn24zGNQrTJ/Ajmgv1I1/gKy8lrXtHa2h1FYoPhqIe3qWEI3SLrcPt31s1rvvXINzd
r/RfxEJ6embpX7wopqIB9kZNi4YkZYM624F+JEjkxmmM0NUrNLaaMa1EEssNeEII32TLDWbfEqWL
DfN7doSqNOZMY0lWgM9+0J3c7OOqvAqWWDI0p0OXwkC8BtTlUqhqH7sTEoYiMHukHaQ8fjlX0tVN
UxiH2jLdb1oVW2SmIVoUvPz6MsUVFxJoiYOm+h674CCMkrvtsffYVMOuXFeOTq6iZbNsMkzLqFEg
iSxzO33jr8Nl8ke+AT35erUUYIG7kLaJFPQvyibiG2FQ3YrxuxZhvPnPILbEyXi2NoVmaaeO5Y7o
wa4aFrRI4vlDYt7J4kBtCQpra9opBiSxuQje0P+2+hNz0NplI6PBEqmpjqLPlKe5qJjz9mCa/OM4
56ob5BIt9Z3sHQnTuUnobQVN8PTXAE6UQMI/4NY/qQ68TlD1L/JAj+43ffMNmBT4rX52eu9BczAA
CBal2JTeelNkr5Bh0TX2XYaa+14k77Afz1LGo4MnEY62CICJYa5n00AUFo/IA1CMNIpEwXHCIvr4
MjVcLlmXjEJyz3x3GUev31GPE6sUKB7gGHvsWR183ZeQpiMg08YzlUteYQ5VfBlYeORekxGuG38n
NuT11MGkifM2q9lMW35aDz4zDDVbChJByulmh4yqp0KQS7tRVsymXRsH0X3vkwLBUj3Ph38bvPbM
jAI8VSaFhAEJHsFWblS/5fRymr4iUZmJ0piySHEz25Yn1rrtLqnmrCNLUhyL2HySEprFkTnAUi4i
Ulfic2/67Qnehcu4gWPBxb06FPTu0wIBxlYsB9khTeWBEnrGTFXCJAh5XyeJEZkxDuRdycC+zWpI
3/BF2CzF5mMYoSpGVvLn6fz68NNsd0vWcOLxo5+ariw5XmNb1G+Oe9G1fWMacxGHGR7hdgcTpKhd
/zuLh6/sADwtXB+Xl73W9+cFttd8LvW6DrpuznIoI972NE3RUbdOK/QjS7QZyLaqrfvd3n5zCuJS
+kce4lxRHzqfy62GHojHg0W/GZrbDIMC8XVbo6ciC7WwdtHbt3nw5y3+Whwhwzu731TDOxEWhBtY
9Bev1V4uDcP4IYSiabgtWB6b8B/liZ3khetEb9V0txOTpC+OvNmZGVtRPpP2v9hxErpHOSDaYanO
b+goWjCxR4CYHh13kqONzM5j9Lu78sG+01L52EngHcCCXITh2PxPsSMe4QUPLr1KNOA40eCuok2T
LItCGTSsFgkRoj8FJnmi68YUcXdc3E3G50sr+t/+Kze4QsWaaUww7GfvIW9B+8sCWtMCJ7RyovSd
gE8wTDOSzgfKWrYtXaeyxCDhVTB0Pnmbi0SZxr9daDRQ9vqpGyxRkgx7nW7qlSVRwYac3on72pLT
HJUc8fpCJ6dlaxL1oeeMfHpmwMg6CFUR3Dde/sjf+XToT1UkKGraJkqJA2MG//81SXZlyypG9MPP
SFO1iyGzv94Jf/Y5kW+IEs4tGfVpjPddrqQ+c2Ri8NX7smym5PDD6CyaupDqGieKOHL0Og+h45SC
KwEQKyNztH+iw22W570QroLSt3nCHp035iNevPsX5uA/IzvAqthpQIv5Q7E3GbWpCk3yxHfFJ2t5
KMJVghsl0LBvFbhaQBNqW4WrDFiuXLI9Qafhtpx4SeagVF6aDTugMwD3QRg8Kfjo9yyGdVMUiHA3
zp74vAx4/NQCsyd8P3AeHCaaNxfr4/SbzFORPR/fVNSw/hW5v/wdK4iVRSNAVL26IJ30TDnPjBUv
CkehMMiVAn1wJrVSqPEGYCUeFc0rnPy02jRiDBIVUeMnrQozYtq49sRqQBCl+abo6PCt3fRqgxA2
QHGtnWHRGvYQ1cZR10WY09utCmIHOCM0np1UVxryhgjPpC1cCPqhxo1tr8Ld/0VtxxyOmgIA9ojA
GAKcC6zXhOmpygNlplvNzGsD1oJvIkTz0GZ7IiOujshtvcqoN8zJe1uvKpHLHWTsQ19/1l7a03+d
xy9JoXW+r9/r9PpOQsV/MwO11mcMvRrHqJoiW1SYXUrX6jSBy1GIt/sWsT2CLig4YkpDetAvW47h
5niTL5+arAzEBRTzybp04VzTKN3aJGYoO++G26lxXL0aInUmZoSGru7qvyb+bicy88xZFTGAn0KC
lUR1d50z5Dfd/c35HoTvVeErW5O5/89mc52DcJ9JcTtKFHwbQcRVNDqU2Pjie54uuTft1+37qrJ2
LXN347yCH5zNLsPKt7ppCB+uwZUE8+RLKCEij6PtD0LgHe3IDouJmZ0yOHvY/y0voCx9LpXXGdco
TKLu5k2H++sAdfR2w5+8Frgk8F1jf31RUokWNXlu32yCQMXSfOAJHFMMVNaOkHBj8nxjO9V6W2+O
t07d2XVEHUJ2xh3bsXJW1nhmJX2grhQbamQNeVZ5tif2lvRMfXCx6YAemQ2Gy+oft74wQcqXI6uJ
K2B8fV+xvrrdbOL46ckrHa9krRcvQnMu441DW4NZtDIJ/cU/Q419LeZSlS8HX0BwM6sJwLWouo9i
PiimSkkunDMZ6kyUfUfolFqCIMy8e4UAzoRpIS10xweq5TZyD2KwnETC84TdE+BDY37xXBkHlDjz
hJYet6fY3JE/kxrrjMBCxImhdTeCv0mR1/WAjOwvIHgemIzQ+vny2dHWY/xSQx+QNJvMeRRD8KKQ
ebeI1W6e6rRVvcHGVvEKBcL65aB0j7aW7/r+01a53+5yko9IrKY049AaNQHjsni/P1xGzz63N1nb
r72VKxfDixGw/S9kfzZLaA9PfP4vO1UXSgDB5ilEw1o5yJ2Er7GxxXBgxIkTxKWMRpDPJRtiTePU
ruAdbcer9+Y9U/WEVhYJ5IB3sosFc8Um5EKJJKquUiF69B0ebyEwNXUYcF6TLW+31jClAhwkpv/4
9zqor8+16xrKZG2MtjCqUik5u99HB5dQkCHANBlBtgBs+/fexZIogixr7/sCdUeaw7wxtESgrAJm
puVOXEEy95yq7ZTlcIs7bTC8xBIZeutYtJM8X8kU6m28gDTgTC2LbmtOfdgm+6MPo3oBPuqrp+Cp
D+9XARtuosnzWeOLxuHLJJA2uCSx68j7b0Qc2DRChY3DISwbYarJpeI/sjtMcU2CfOh3LLCcii9/
1NiiP7hkHWYmsc6l5qau1yZdms8Mf90UjGLHz6gKOlPzVXzyP5A6Sn1tq//1e5XSHaVOReJu/OrV
imhaBvlzQD8lu3FTz0L9GJzXSQEVk/jnXvXieqScdS5495YID84VN/QvMxSR8ePa9p/2XRFjTO2p
bnfDuW0ccOud56Icw5NORlCt631Y7q4NENu1YV6WJam6eaBgYWFUp2Yz66CVVpyjAAAp6ijTfDoE
rOu50rDJhXCu535CRZu3049Xmcf/k8R2NuQcgQj2U1cEz93EOEvJ0yhN0yP/zxxyb0TjTzemPzqh
185ulDTQ0KHr2v+v6XAabrxhglxcO3wu0NBDOENpHnt0/1DFOLVIn1UOb5ffVZILsOQX4TstUyPs
iCJI9WHkSqLetrQEV1Ld7x6FlejGll8NXRnow7AARMPxL1qGyfdJPA60XCKQ1mZIhbR6K+n7MaWH
pvST2CYncDFcWnd1fYQexBzvvw9xIstM0ecj46DILBgRNzkox1BRSIv4zcmjBz5RH6xfU5lm8C/g
bbXcevsZ5vg53sT4MdbNG73Jy7B2eYHW//YM6SNMxe42OD9VnOq7SOVRPmqgYY8Zx9CBEXufDaWx
W1p/iSth0lV4je2MIreXaX5mkCKdHzlP5Y0aMuI+PevyYlYT5WnKA2nXZDNqt6aE9ZKu/LHgZw9m
g25ygwIh+T3NDWvAbDzaUbNfhkCAZ8oz5lDwO5o12XiUjBXR0udAhMwwxhkijP4L/tAUh8UAzblw
lkGxrpvVjLHOO30HW/4w0F0iBh+Bd1qSzLUIovkNnth6bvjxOf6Ae1nzYf8D+6eLwbLT+eKEu9vy
ZQq8McoYZz4WY6ZzqQ+8TUzcGMl2+p6x+w7mltNTdSfpKtdPc3yFhLHbtgS+HhqOaHWbDK0YrRDH
o9mbiSCU307qm1pDyyaBr46qhvceMUVghsU6+kbAFt2GVkppPW1pg3kCLQJvL6HDKuGP1Muipwmh
53BaaA3uz6L7BcJqX5R9sHYKF1wC7ZHccZM95XwSpNi4kPaqWuOt/7RAw4tIdOZ5wOAMfBlutgNT
rqTgwGmBidVUnV2MxnbDwp+iobSPmPxl4/gH2PD6ta29pz6I3kr3y1ya3eUNvwd0S6K0WcOAsv6/
JrymECW0uWxD7Kc6UFqgZUrM5cLhSWRp55wTJ1uOke5yEcFAXcH9OEFlYvDczmDogMeBHVuIdVPH
jy+oFbzZzHXR40ufwsb1MkH2XFj2+T5UHipfmCxESdxFZWoCowyou4lXs3EDAHhN7EIPgLEVxrKG
ORZr7tUYFyZQJv+kB14QHY6qNfbuQVHpdIaxC1uwTfgk6Zq6Tb0jSQNQWwzbZZyZ/jN5H+zgCjLD
XK6HBP6sSyljZJrdzDpdGdplJAu5IyR2MboJC6khphy7PWkLT1CsLRhFqVRO5bg89SKH+D5JAZsb
l1RFehV/LEKuaaTJXGZoVQLy9w+evkZRlmrDVbevCYe4uVZgbFaCaDItrvXD8KapyIDF+bEKsXOO
YicDyQsaoR3XGjnqxJmanY6bMAh+KhmuFIh40x3R1O8ne+dpVSqmEumTvpyOXccGeLOcOMc52edA
lhjeeSLs4hzeN86WBqkC/4QewjNaxXA310YkrfLs6AalrjDU6jK6FUhvpj3hSchCwTI15dFn9Xtj
z00I6EkJkZfmM2JQVr5g/z8E4juBstg9yET0oZHROBSY2FFJMaVCmp56C8g4XuCVI6vinSFcHZfA
FgmcpmyoBoGzw1UyVzuSlhbcWz1HwHNM4/N/uTFAnj0Lsp8Qz2+J8nHIQxAcfcn0UyRlfFjSsGob
RcQnMaq6Dsc+76Kyp5ZsJaBznizLEsbxRkKccDKDgBx0gS+uGJ1C2rYio6WRYZAtY+OvVNjSGlAU
TsXahxYpcSRfwl3DcBvsJEfz1SKCUPBPBT0d+u5FpEPuyPg201ezamCK4dYKtym73Vm1irOcblyA
Vos/xn6lGEnx81OKN2mLJjImA7+SQWbDWgNPU6VzxAbL2d0UF4+W5EnRXYAX8+tZeSt1+XMnfzD2
roSaDOP4UoQnTNRCHYhEYZ2KT8kk6AOorivE/B9PioP7VFm7n639CzKpO02CW1S30lH770ZN9kTr
5xXCiXbIx1UUBjhVR+e0GwREWI6v4BHHjjkjeQUok0oqigfo1ZIiGj4DvTyOl+/FO/NwzGidVFrY
eOvdq3N03B9DeJGIgtJp7PZbOM1TinrWbDukHOmrEAj+lbWRYJUfAeeuYsB6ZKoFB1LG5mlOMi/6
ri853Qq9IInownfj05WyZ99q3ydj9iAfTrkX7unnD45saAuHdfuoZWKIljBwb0z+LFnvebJOUmSR
tnRr0SHSgCjUB0TDSdFl0GAjgeUit+MjhKxjPA9Hil0IP2NrvA+VuxFhfBI6uagq6mYMwhbss2Wc
wNNH3exAn29j+zYa6YGhz6JguByW1lvm/5oGmwhlWfig0ivYOQ4ZH7i0c3526KbjoMdGmIeeDVJV
O7+XfBwiSnKZJ0Xw/rZZMj4U0GPKvfMYOVCMp0J2BgFkf8fL8QnBXGtVuUX1K7N21toBmRbBVljH
uqh2jelAd2CyMAZWPqtiFqEK+PP3c0tr6++Hm9WnGidyb0RB0gM6PdGbAg36cL4ULlvey6/cvExG
93w1Wug3YtU6DtuEvqNo9Fg6n7mC+qpBuvXQmpwgnYLjduyOX4ecNcz7Al3EGtE5QzCghYdvr4Hb
TBKFT6LUoqVb0SSAdgEbzc8OuwaHlPut0vrDUwcnvknK8LGcuskclAOMVmxq7eLschHwtoQiUn3L
bb+QaWAQeV9KTMuH+apEnTzo2jcZa/pvOFPniko5jzYpjTzU8qotBuy4r+BY6LwhYL1+A/EjIxSa
f02WQOvfb5KfJVsPiWu7ENXR4a+7nSVrJWnkz8mUw2zquKEVAjEg03XrDoQtUMiY2QnhwX13WMX/
2RwFb2YFTuA7AU2EH9r1Tdz5fQDRmPYAeZdE4hOLaIyTlj4nzhuWyEjX+J/V1mWd0p2BKgzu7lja
fBh9Nb0rjhYOQ/hxnAzKBlhprNhAy5Ge39VBQTYtUk5DDftXq+wktyklQmkLlmOYTmflOEB4e2Of
D1oTGUXWNKNIqz4MFW5EOywHi65+4u8tu+hixfkOdICXXKvy91tDDhh7/6r5KAwtN3N2RKsNGGUB
VSqEnOoPj1Ilh9bhN3LiK/nGrulUeMWeAvwlNYmCxc8Sf7UqmmRCAe+8v35H68ephppIwkgOGYHA
S3RuO9hsu4nBbAqCHAkbiWX9oTFtQZRNJndTY4ffBkmmeYL4wKiQbBgo2kBx9nqIf9CNE+dbTCk6
7ZbtKNCkEqMJB6OqgUP5k6pidKdA9BIztxTnfT4Mp7KpL/Ykdc7/benSNADrqG15a1IC8H5E/557
ygxOxR7qS/eZ6W197SvinBq4CmGPEQRap+ggfWn4erZ+UIrZKboA2vD3Nka8oq0jNC/TsjwH6ES4
3Buo+rShqCz2sFsES6hbwWOnn7vzbUBNO6AQYZdCZYWP5tctxlZInZD0e3a9RjeIF2b0Qfbf306U
JF4sA0tEfIlHefDJhoIC0aEtM0oMsuOG5cKK/kIXerdOAHNpd73tMemFzX1aPz7z04C4WZsFpw5m
pQFoh9VUjzBJ6ilJqHbLa2ay906txcGhl/GpqofU2f7xhR7hko2+Fatir3kSeA52lXsFtC/tbkxr
TeJReUrX6GXjA1VWpZsZg0GjnocXndtu8+Q35WIdDWaU99wxD9W3wnK1ybPD4L6SxBlhfE0tH7wC
m66tAoiEp6hvJW+ayrj+ruIBzMhl8XDZ8jdMdspJmbXMRSgkfIpgElyyqSaNpuOOMLdsyi/GAURV
pfkaW6nh3TkqFxnj3hx9X1Opq48jF+b4LsMGWHix/BH2SLbKog7jiL6yI6MPzveGwAjkj+DqHGuM
kmWBzWoTAGDBarLVM9TrXkobozj1MYeLVcqS8qpPa25IiGbMoMidxgTwFyxUFwIWKtpjZQ/6XFOC
b5NRdnc3MoOxbthJLfMCQKiwxxhENplK3nZWRBkUOXP7Csn1iaudQgIKd0llpqzA2OTz67N+jlB4
biT1ULiPdFr2YoQ6QxfXtQOx+O2Km8mGkIzz6jEOP/nqT8XurVX4FC4VbcTVPwWqYRrf/Szb0lNo
4A5XUV3y6i2rTqfGniNODe2HMs0qfDVjeMPK8guNEa2DoNaRuU6EbqjYTgGjVSlZS3Nc7StssNAT
BdeYClrfmDkJsFiGiGyqZirzE/2uoFN16PwIMBR+xJWC1kSWeS7tzIEV+Hlw8FIDQZ/7UHa78vWe
1nEDAAgNeLeFn3rzpNmGtyhtQkRXwEbFcDOo5pbot1FIbKVIrUgSwnzAj/AE/IvLZitiYCmlbECY
04+jgjMG62buCjuhmAZ//k24AMJ+ueuhR2DXtPx2gyHx2RuNN1j0UF0/m/YrNVx1ZffNJk8dKUuE
xseNtsSPLkNM2b8TXjLoVl5JeDG1tspdRIYRIll8XgS9FEdX4AregdZRuh887NNZHXKQB8Qbky6A
Nee5szPYIjgl7d2rWpcfkPnepFuC6a99fBcTuwXcZSlT2N3N1T1GbmeCiz6nnI+leoQiffoOQ2a+
j/AZimtfVrYKL4PIiifSBT2DNe6OA/6oRdn4ywwDmMaaMa25qHXq268phKQ6H5Q6LvuzrdporUJH
k/0NOI50ilLp5+qSWXwyx5IvXq8APzB63O2cUdNoGqtOO8dRDaDBoOiP6MqGC0GnnV1Piu8IGqgE
tctGL91srOMbd7gnk1s2SbsTusYQCAYiEYVaTnTWGA+907vlXvGP0ahWdTSTrtLGytBNUfx9TmzE
B8qqpp2gBQCnObcBMeAqgmk6rBzQHfkNXoq5qwKttLLm8SAcQoptu2NB5z0vCN5illaIlZ4SfMdl
3zOnyzgBxK/6qUpkimYZLPVIXSHmXFi9/xaWdvyIJWJHUScnXkJIAFeYM6JI86YD0KPGRnmIM49r
oDgM75BDcK6v5lj1EFER6Zm1+c8z0/XaR+qriN6yc+p3GP5Ha3YNMtjI9L9MfpdrYxiTxNYWvi7b
6XPBzwi2ujoyD3sAAI0Rxb4JhbvZIKibBzMUOUVtT5Tngei4f3vqe+H/OTLHKKlDZdsK1hViar3m
XlVt4/j4/B97NgkXduo++e/dQamn6J0gAd0hgDpYNlG3sbVdE7x5Vnnv4KJH1yK4nuQNQrrIlsxC
bcRaTdRp2RPEYDzCkNWk55JHYZXpcUXmXE4RVxgR53KoYqWbokokRDhPDW8sR+s3tRJb3oaJa+ji
+lYqeVrITiuikfrostYDGiysDkuYjpnjemijysfLo/yKUZLBdX75xLcMquB1kq+W/FlUCUymjgQ1
NK7JAE0WP8xOFyg12fQ9sfIWXva+P49pLctxdpW5xCR6r4Jr9LrHpb0zW40Jvy+cUx3UAP1SgUfd
AP0CjaBHs3R74T19tPjkl/J1Wne6/5OnXT+nNxnlsHJMnVObq3gp9Z6gvjwgRh+73nnBpfCab6gF
43Qa9hzmW/41bovEc3yiCRV9FNkQXViq09rhe9K3AlhOdHlR7IapoqJML/SalAYPjWDiJmSm3rKM
8S4VOgj11c9SEiRdI1I8VnE5Qaq62v0Bn4dmXrd74zMcI/YGbkN2XABYw3zbvMcO4lVvJdJFOp3a
RlnGFAflzxavphWYNzuVCzyAfOwSCpZRshY66YZBynxZdZ2ktUpxbztTKjO6jRZUhr0qYyh6w8Y7
WP6MXjUKGCuYa7h5KYFaA4y7qbmJazOpVhaGo86Gcz9uAVjqyXRHcVyVPmXOXSfVjR2B5IKON1NC
uIlErVTo7d9DFoNMg9ujFwULJabJVk1t4GqNNevkOBSdAwreae8q2dOil8vHqzRkuB8hexspbnsH
U74F6xqlVJvsQSkgvlQHRZs8PT4aZFwNsohV7mXMimvI8klKTk3rjNnaZLRJ2ZyGblkvCCPtCvB+
l3G9ZjyA9vavxPixcZukTDxQ58zYBJQJrgpwwz9RmyRA+DB5WdnOd3N5w4aUDiApUuD8hwRXcl4t
EH7Tb+Zn3TMkLHsnHlUIcSS9M8VHVcFQYtSeKrzPHU/3D4hbelNNFeyDCRIGLQSLKGUjR9AQnQcC
ZJi92WQc7LMY1nR/T8YhZ6skw54XbmHlxvFotrxjPq9WhNbGTih4o+mtlq1wDiRQ+28JbX9t+M/m
mC3PXBjTPzwMgrSLQLj8JzanMyLtUhKhc2mzuLckbGs6z/uKXT7qHpprYDRmD3dq6joT78/PTUdk
xElECHcZawEVcDn6pCBYlRAcceBk4M2BWUfBgDtoxi2Or3CGajQoBxTvzqjtA28uOj0LGOCz6A1F
5Oqm8dzB1CD1hI5YoQPYwRqqbRKz9rFoeymbG+TkuU0ayANONpizKzhfUkpac7DrFVYHqPTBBepg
rCQwZv9Km4xmcL69a8BdCNbScV/wwR0EBFR66J8GxRx2NTGUrXXIm0l0ZrnHx8lcTBKks/1voUnf
BurGULMqCRH4y6Hrh2cxYFPE3Dc7YV7rKSqTKAQkhIWFjl7JspvdJtZUDW+5ozm7X+a4zYFWd+YG
mIOGkGx36lqV9yfhTFIdlHsfe/TcGRgUgdSxxC8ORKWYhxe+7MERe6q5XXfhQKZO2o2V17mnfpxI
LhydG9HJxfpKmiyeH/v4JLJxvF3tNSaR3lm1baYf3iHGhx7+p0E0LwMZ2bUw/iqOmMGz9kz8We24
E9qF8bQ4V6L6q8q36rtWv4D0kYYedmbaHVCJWuTFJ438KEVeDxhoHnc9LhhAhRg6/1+dIuSnbv/3
QMtl5o6HY4FVAmqcMmeHmLRZbjqx7IuG6PWNC5pyzwZfOcPa6GDzRfj/seyZhRmxylXTWOduhpTT
PIVZDQN3edQmN9rR3z8mv1tJYOrxzEu/gkIOtrx1acsXeXd1Ewzsvpg/MN57S7AEJ2EY16gQ29/D
weA4hWB8qlPI96L+B1jWyBzc39K/CSB1belDMwssl6w1Bcx1y931xxPOFvS5ETKD9dcffgX9Q2Y2
nLWBi9EF2yau8m+Dk8QdLhWrD5XBbmyk3PKWhJn/B73BiRR45HNTY2G7IA4NyOuOjmxHk7fsiGjp
fyfEj1vve8Ve/QdMGr+k1Ojt7dbhKgnrHovN1USghxMdwPMui8rJgqlFCVJD7fuZb/Rc4GUyva5l
y3+xclSC+uPb75NSg75rcrNaOChw1/Aoiu5GM3vBHE+vQcyEqDlG7qWmTfTiUNoCZvNG8F/TaT6/
1aZ8/P7n+v1sOLLt9u28XglbVDVfk8mlEwFirJv1Au0Wmsii2h3fYG3OJ0nbTnfUBhy77y3RQitD
cNxuNIpAnOfRV15v696tkLZO7ibLx1bNcUCiD3Ogj6zkCRngmRDxMCHhXM6bZICPCkrDDrIYdgK3
zuV7YaYLZfPU1ykO1sanaWSsJuzVe+MsQ/rVSQB65KV0zrJTH7XhY90vzCrCRaKd42ZH8sbtqzkV
nt7VQtUiMm8nsrfpt1FmP30uYFyxM7iAbjklUyTaqSa9AlB0INFa6cJXw7UPIKWWGNCAGjHiiLuy
B0+hnL++ifwzq8nhX76/REtqupqXiE3VXLhf0uY/4bnx5H+y1ZeMRELItv/riJ7rpqTb8Pho5s+7
YoyPpTBWYojQvl7i6wFnBLef/px+RQclziLzzrp2GSK0aAcDHY+3mDuXyfP/6Ly5pJB+rflj08km
kivzslebBgW08884zfdGOpO4nPwcddx2XgovBbT50KEzaP0AI2O8bAJULNGlJp566L7lSwDH0lk3
SlBMV/t1CNanJ0uGxChnz12hSqv93h0Ji0BBQfQemxjiWfuF8Gu78RVGFf3TRVtLE0eVR0EjvJZt
Oib6yEjSdVqAdCfUnptawzgT049GfkG/BMNIh2HdDA+BSimql6RKFn7LH87Hojga3+mU9rD3zkPh
tyj/8zFYEZabstsk2GXsUTHvN8Jb/rSewerfblwP9ekzvvHOardLSjCyLU1om/rjONIMcz+bfzUA
GEHr3fKKhtsLgYIyA7FDA/ABRG1JhkD//Xs1yG8dqqWwfXqU3+zhG6Qazx7CSPfaqSL5x69BHvzD
LAjzZg/i9PGF8xXlucVPqm82mucc776rTgTHCmmIFwGY5EROmlXvBuiXZhNiXDALyckZRaq1s/Ik
n0i0VHdCvOVh/REKTtvw5aFq21kQkeFD8/EyRGefZej5JsOG1AejdpDqXE4+nuApqndpraW9xO6H
S2R63LTP0shbS1fo9kniVcbVTa1NjO9dafBFP1tN6jAoDNh8tBHaw5Tu559wXBPYzQwGDsTt14cp
WfAewN1T+TUZbwE0Ku+7MOe3jEAPY2tEV9f8BwlCD/0HEc2Pmuxg9NFgnWZoyazlha33DsJKRkjq
B10OKu/8KDczYbC+MxAxU4uk5SF3jxeK0lKjAZSwhnv57XLr2uRm401SB9eQHZcN31PPJFE29i67
xYHDOQgq74/WtgRmWnfASZZE76FY0gKl5CrXvRUihjbOisilr7CZX7iE1KeCNl991bWuQnP1lHp4
dSRmHQUmTiMaJJ2IiTLlVgAdwIALV3fGyfT5n/cO9VjT1FojqCk8AK3J9hpC+q033BKEBK5bMqlR
qfCxOToQo5KYuhpobeDQCYlCNrSnQ6AIOBr49YEmEC7CmgZKKehKJkbNFD8rTRGoMKFI6PJDjWrZ
MCcXQPZNn68PlwQ+UpMQwJTXP7NBPbUVTQa2dUKqJrdjsxEekIzies0MDqpxxPVHx6kwz26YTV0m
CVifq/fFxb14et9RTjpxpqOLtnYVxMK9QBAdc14xpF8Na8t4SSS4T0fB2B5aW6Pa9vNBxJeWkNbO
CVxPWIdQ0AR9CZAbBd7RoSNnd3c51E9/YBCyYggUJ6dapN3VB2lf5NDxG4LqPWmJZH3m+/3rIQbE
rKwIcLC8GCbiGPiP/Ho9JFtiRloJ/EN4bV40xPmM5mk2SZt9gAekPbLZLjEI5oP+67KgG3X0y6XB
/uYppdFssfv8W4VlJBioVT4NfBmMtftDc+j963I0avwUapPu6aKzg3KlYprYMHNqbdjzYMcXKxiR
nnv0bZulbOW1iTeY/Qbvny5OnEQKxiGuLwKV1RKUikd+9AyO2+z7R4+y6sGdBrujwHRyGJv0F5iD
zeK22WoDAiZtlMlMr3u3fMx6He599BseW28hd9K1dth4a+1DIUAS79tB7zSfqjaHvMz8dOyKNH9l
8N5VQi7oJNfHZbq2KmnzBeqfdStCGypkR9vBZdERvY+4aT4ctTUK2aqKgj28Fztki8/lMVgGjIna
OPA6k5HuzhkAX1PjldUcCd4sN4gOkY7X8NzRakzOtFjbOuVC4tOtypEWaTM6QEWT7fSkmbPzRQv2
C2B0e+S+WHxRCYbUOH4RC+J/akvRt9UuD3YF9ABhT6gHGJIEPEc5pASYKSEzdiaCLZhVXJYLANHN
HEXjysYHXHhFqvjFDCd0CqVdFAtUN1cGRl+ZieCm8yqgsCSHmfYEKJs0X6itNsOfGQY32VDvKt0C
NfTYsMpmu++6L0szmRbYua0ri+5i26meHpHVT93lEnSLk8C3fTLCzLZRgffTb+X6WkhP768kf6GY
viKG+bpyeq6CI856eaifelZFdeOME5UTtEE2zO/kdxPqcb8uJWajofpMmhOvHiq4Gzd2Rw6bE/vv
bixfWmbcUU6OvtjZQlTSNa43ngrPFY6arb7V6N1E5b+xsDYpUmUuGK+/61sjTcO7i0lPg9EnchKi
598fDrGaIvFaY6Nu4HBTO7qCODOu1kJgKiztkeFp+GgkJYesutUw6IJE8QUKB5oy775vWazjVPuB
yjzT0nHup4NkWhcNu5/XZjluaOjNYR2MYV5zKXzZWkxNC45P3vbWxEhOMylQTwU72vdpIBs3FjeM
dofXIYGogxMpvgT5n9zH8jefK5GMt97n4ePyw9CbRVYK9UPUcfPLJueKT4LU5GqOVhoIBmRuVNKT
yfTMjR/ayv6kwlgIzq3VNjcRkXh+8ECb7WL9+8xzWY/9FNmAk77nNovOk2bDoOZcR2oVMpMHL/C9
yoTWFVCaRigNgn2LdKaYLCc7yCS5p+enJ+/KUWFG3MT6LKqHZZQK1Go8oOlR2azPOcHVc16ColxO
HFe5p6cR5/Dig2hdjoOg34xtx+8QUgzDJGQfzDcbLYElSpdIq5QSacdag5ED7Bi1Wtlmq6Xw6zza
ixjsEtMERhpywIxMDipKb2DhKeSXxUALymwDJMPZxWYr59i6zl/f0XqEkQgmlNBRHPSE9iWiU3qh
eEw6MDZcZo/zeNeNql2ji/EqZtoi33KxMiPG51+fEHMhU9WBTSGevebhiSxXs60adGbYk7Y8aEcT
BU3BerY5CbdUXHH0xb1aJneHub4mFEGiMkH9Czd8hKcYWjxcRcrBNWfzyHYVAIjKRrdiM9LBA2RT
dEp0uzhekEHufrw3vr7i5e8LZHR5ukqrL/nVWsjrQUQD0D56jS6P8L3Tq0U7RNitDhO4AsnKEyDN
x4D66+4H92dCOCfApbRGwPTlx9038hT3xV+MSmBaxQmuxTuc497zZ/BOV4fwjnYy6MrItcI18MyJ
RHLt0aitsyGgQSAyoSnzgINYd/3sESNFBARKkTYV+YJsZLK0oW+37PaKM7sAyG2WjYEUERSrUIgD
CzmEAJ2RRJMa9HVWKepE1wYnMqzSNI1FkQ6ErCwyHQ3ECDBmFoRIXrLMcS2FrMZ/kTmLdfvlzSam
POcZhQqoWA3StglAC8geUJBrSpdaOgJwYeIaVF6h9QXvUcQDNP1F9SwFJyKOgJZT2OYcaSrombA2
MKeDaJCfLAa96t0mzd8lAb2WrKLbWA8izfXI1DHZICjCvVoNruFIqTneJa3H8SJt+3mHy3Q9RmwF
IcaDFEABPruLjJRu/eOEAjqPXuZ1wDRb7xjTjkExe7B4DXiAtaccU4T1ttPL6yuD7if5gxsn6mbK
bbVXzcRtOIaXnvQy2BtIMgsG4DAvc2Ic3VJmLW/hV6OmZlLKYTrkBHHzEuZ0WxCgZGz8xunO26t9
qvk9brOJXzyG7AFd8AuCDxBA3/QWDvuS9mt345nCcaOYjEKoiCjC3D1wSZSN5BJC6J0S8yBdkqaq
iBCvzV4XsjUAM4ckGIXFIkpNlefdRxFZNOAIwuosAk25i3t+QBbSrMwkp43CG+ZuMu1D/La3mo0h
IXqfzK19mN+KLu/CqMY+9RpEXvMNH2MRdG3p/4DAaPM5YBQu9byLqiBDB1CohNClyPnsjmGPw5J5
iT3/WrSeb+h5++BDr1pwLyapaLngnvA/pyhuYSWQDIP8rjEB05c3hdGvc+1dpO0rAoO/93Vlqc2x
/wqNg92yvVX/FIi/snyRWW33ophmabspkoM+FN+X8J4uS7DyDKkazbEZbV8i1XLfRKSh+38YsUfE
4MsLF/cREbGtjLll4EOihNosE+Inr1jDrEKdrg/sjvBiTYjy0BQLjxfg2S8Yi1wcxiX8nW3ekUxk
2O5QTAnFcGbwujN/xKfpaZo9IL4BZs2vsNjQRGboSBxicQuh/XFWqWSk5w4o+0rXdqa8KFXWfP+o
ew+ttr7qZRYM6QhwwS7NcU16VhIhgDf72Zo5bzGRVW5vdwe63c8rZ4uKpDI1wDozmOQ2UU0cagI0
Jh4IL+SQl9rkKX04d79+vgywXc2NKzZ/cX76yEPBamZtHpYsFKy+R1RZSvFf+jbsAXFrSyH3PN34
VEtXwKs9uHuYQkM6hyO/Ld8s1YCNQQhWEGRpmkFyvWsPNJw9i5xuaPa7OBsjL7Ecf5yJbAQ8Z0hl
pBDfA9WoDH7RFEOGey3QI1SBO4GupCczlWh55QYx7hgHQOUe6pd7YffLv304T+Rjn36d+NBztO13
Ob+f7tDcTA8rXO3BT7zyEAH5qcLO8PQPyxZ6FkFfNiZkyrpaFkDVa7bI6v3nZyv7v8Q513WL7+kQ
b65fonSEWzytS3lv/gul0GBQOWX2u+r8LFSTAJfkrsJzFvqY9joaA3i4Q9n22jiUBqZA5QUVoVMe
kuepUgzSRF71N+eMtBay18wtoL1DrE2uTrO1wkIDKGCpjLDvzTm30+LiHJ/HQeVv0b7tnSvUDNXg
Ow8ps/WYlgZ57cwBJF5atuzHGJIfO0gk0Bd62yNXHSYV1uppv8c6cq+RSBHUbSl7Um4bk+EFFIQf
NyTj3ABhUB+gPCEz4shl+PbO+HTcuzyMU6YhVrbuEDo9eSV8Lw5T1mrrbBWe1rrKRA9OowZEFLik
IJ+61RGvgEjo2pU+0JzEOxNIl2W0o68+nmde6ePMwog6HPME+n67beb9eCmkEBjf/oVKh/20Ei+I
nZvW6j+LFueMaXqf/YyndLWhQMYLgwXSBxlk/ne4PKRBO4s3OQJmT09uOloMgGppjbfQOhrOfwNY
5nhMDWFBYcA5zZc8GMWhsdFL9fuhgN+WLUwb9sE9yH9aiJq2scswn20ju172DhCR4e4dkKs9iVgi
wn28IMzAdeT0AH86Bg7znIl6Ye32KJ4t5Nz2VqrPEYzPRoJeMpbVDU/WzjefGvpLjOjwnmrJl9qT
3qXqETVbQBt3bKPK6JnlTu5rbN1k29K1W+qvLzks4Uwx7PWofqY5WjeS2U0QWah8p38YOLGJydLg
iPGMnssaNLm/VLMc/gEn7Wf+e3t3tvlGMLePFq5qoBOWbayqllYjAME6C+enErIUBkCbfk+9fb98
QiwueSGnUSKMUQPozQdwcgR+stepi4uowD80d46AlhS1Afmu5xh6tya13RDkvYeskpUTYlIwyxP1
zW2t0JZVajIaEcc1ZH+wa1gvNxQgh6Esp2F1VT387PT5xgEMSyNYRFLZbKf72+qpw5t6KeJ0rChU
ibwXAripKUjRsZDn0bg1V5qGysW+xoimpws3uMI7OWSVBM35jD0VsJIUXLKsgVzsF2YQ5fD2Mnac
nqR0pIPiZZ/pUAj5VW7iwZDiiwC4sWG1mRE73bCbpzsJejcHXC5/1VnTSLhqFafgR0LUlYNRu5+1
D8sq5NKkKMEzWdm9hB/0R5qN465P/kz3cWwi+noKgaTNHN14C1omibMFJXeaheGJRqpapkSLoobF
BugzY3pZtL3KQZs9rS9IDN6eHlMRpwHqLvjzSCQAWiShtd5XWuJ6ZIfwcUjL+73SEUSXAzkxpai9
EvdYNMZaYdhTO3/8KjM2h/tUDUGE1M/PEH0fpwdvRRskJ56ZMxNsQRMn40OrwcgqsEIfkwqfPVO/
YgZJ9/+WbQxM+IvBXwaNg7iSuKhjH042V4tS7A59XPHHRhhWbWK1W5/XSbzNby3B8n2FKTNcMULu
S7BAhQ7ITFT9L0eUgxSACvaKrqFgr7tFKk2mY26Ait73ZbNdbv+DvYS//Lckykgp7to2x3bQkHIE
2kAXl041rOtQ1SpqOI5GAKz6fzpOWDbSuPDradnYzzPIuf0srn4pfluOQd/G9NiVn36625G8fJbS
LIMPRQE2au1iit4zT6Vj0LzknJ1NuVvDoRdGdUa0+6vAntDyQi8pyDVj3uPwkocGOgl6zBqOgpqd
BM/f5CCcQklnIEBGeQGXzTWQSManMt9Xc+AK6rVj0bCjN+hohLvNNS1Q+r0Ugsy7lYBKPyHVW86w
/rJUfSpn1TuTbx49KlUo6Qb7vj1Ley+YPfB8mi80AWHEHbFxlHBvdikHNzUEVs6vJpNF0QAzZCZp
UCD8mNQNj7KNhYpd7cGU8j0xU3F+uaiyFnvSzuATWDGDi3e59bhCHytA+bxvJ+19fCgDZjbxYFd/
KFfJy7InS/6EOzR5ExpBxUL+8RiMZs0/EsWAOAXH2P7wvF9xSpUw1++HQ0ahDxXmC10Q/Tgqv/4X
M7N3Cx3kjhld62ROdZty4JDtInGGQoXesTWXR0rZ3lv8PZuPoCTmFJNo2spY0XPAPzdwfPrWxUWR
gGhlIqnlp16MFqVyPxUfAx8SusXSV/5bo/ySGaG2rR0r8B51ZgcbNZefdzyCvgwmHl6lj2rXD8+3
GVF9Cfv6933/zm5SLJNgG/t9XqEKoPEWsdXOoC0nvCsATHFvz7quRdPlHN0grncGFjsCE4KkNoR5
UWw1drMJxTfLU24NVAFjvjsQ9I/7fLy7FQV16dc5V+2Imlrnxk7kFjdDeWDgOwfbsU2pgGGO1vHd
43US8kCSigwrWdySvrtkkc9U0VNOQtTTQX+B9mNuxhIC9kPU+k3Woa2nv3KXYrc9or9/qBxQ2cCM
6UYGmUAz1lh5UrH6oa0XTStU4DqjCoAXkunXG792fFMb2tsYZ01/qqZCW+KYC1UHT6w+moaRvLIC
5HruGFwrm/dRXhnFKt4lNKougWy0aBeJ4Uap5dvLtBfv8c1qqg84hWJuEpjUcDBGv8P9pFi0+ZGk
J2YH6eF0WshN1plChKQewkQ7uHflILSiHL13SRYRznfeYzi+xbDU94A78LG1S+hS58LtWzC7639G
wBcKJtZcuxOqgjb0/lgNzs8HGxO81ySf1BeGDNYqEXLtHWlfy82d9wSCr2RySth7J3Zmf2YEgrWm
o2TPgzmNcQ3mn2uA+GjrYP9P7jwJ7aHdxCFF2kFFu5oa+gnFdbd1yL85lXAQv58w0dfpyzMsQgc/
E39NWfXMFQcRnEOODcDEc7cXZKvHIrq10xrutnXQRyyAJ6eH9KT8GY/LF8qz4ILweOO/Z6tEs2ej
CuacoOCohDyJr5NP7rPEujI5HAyi7uw1aoagR+K2D2iR/rLUDSzhHsElI/FwmgqRAYoCUFCUXC5T
M05yooYs/R4DMjKPHMzYWLe4HFoDsjLZkyMC4xsYL+t+5FIz4FPn/7X5oMqu2dYDFGNJJUknLFSL
elzNlcHxF48vesZtU5CIiXW7HWfkJ915RS6QV07zDAX8vjPCTIL64mh4P49E8gNpZL8vNNioQA4C
LEJ7wLunfS6JV9B/Ec+/kV4Kz+ycM3j4Ca3pjbYf1TjdI/o6VgcpVWb2vCg8bGTjyeUCh1zbJSJC
xFduv4+xqXjFD3Spzddgjv+tp//Ppc8p8suV5b+lTgrk1+Yar7x5lTIRcN7wE7UWKHzU8fNLA63w
KFM0BEpwRYmYvGxjh0BFkV8TQu4wLpgosWGivtxZIy+FOo6FRQUh5OlCzqQNSPYaItoZPQ4d+f7m
6ts23Bb8cp4qaXd6/q6ef/DDO5ELZ4CnSsIeOVQ8WHqmflGXGXDCoCcSHZxhr4cgb1jxZk+KPZQN
YJEwV1nVxhY6L/PHvqyBq6GmyusHqPUDRZMF3JBsGGgU+OeQp+6sP7NdDWJegQVnTJeqA/JEqNpM
QE1QUQOcdf5nju6ou2/4bL/YRscw5EufjU+6/1kHxJCwd1edmW6qUpIeE3lBw2aKbh4ugS7csZ0a
dPq+ofrfQqVZ8TkFv24YVTmQ43s4GZqmSt+fLCio80QycR9ZrdTAyK7/0uLz9uMMmpy7d8RNWzDl
ZCHCJnlxWCQFuQSADD8sEtDyk6ZuZrcdrFm05vuUFH30HXBNeFHZCGb2U4OLIbWG7jw9lKaNWNuX
HOYz5PoyZCO6gLyUejcLh/emJ4ahVZOzij1Zukl9AWxs1UtrJJOKlUvLxlfM/V2PeGNPPnI1YF+4
dKyX4DFy+ypwDNnehWHb2cJFaY1OFCDR6/iWjTgG3XCdpLKcgufSA2u+GurJxZPbeNrPml4Cb6QX
uXsR1r14wUy1C16nu3u/SsL+RFP7H4s6k1KJ8okxWXF1jzIRLm96XlXP1DX5Vk4BYdUdGxJDB4fe
qYbGsqROikViBL5DVewV7eqfiRvYC7SOcBwBJre4fpn4D+KpYaEXl0HDy+pgthdmxUvo24IYVQjn
xdBlt50mF166HAJGLty9q5JvNs71+1GwAKXTHk+uibGJogQEGkMfKaapmPeQAvdKRNPOuXMLopHa
8cf2t4WuDmUlRvRKSmWsyAckpJmhyvXXHDcdeyR5LPvFmO1r26iJHxlKirwos3F2ZuSEUUWOX8iK
GG4d9/7FjZTRUhQ4h1kXpiZc8tDZ7xNkz68dXg7K1WbjXA1YAP8tn2LVEgMPcrNLHdYhW4Q3Q55B
pODBeyiUKY2JQuUAq2g36Iqbe9HZAa6w0LWyqvOyrC+4kd0akooB4hk0U4FhPqEm4AZbp8Le2yn8
7elCTZVPKe8ur6kUOO9eGOoco3Oq3Lgog4zs0r/AN+91Brv1VPG/bIBZuI7d9wV4cWSvtxwqK6Sn
Z1uNWkUqeHt1mKPMsa8rUu4e+i4/1xZL3sRMvmxdZ9vVYDEGoS4cjgtdyMkdYKCa1XSy/gnnjPJF
b4l8EwTMxcBHG6exa+L1+lib/W4Cfcp7OwdVXqSttXcKa32liH+a+2N0rNBfeAhNzZXHRfe/iMkO
mPixMNvttCA90SEBiuS1j7lhyayNYi080QpTs2cko/jgVl0qTuZXygbds5h1aDA/RJD1gDFpApNh
pcmlgenJND3x6ey7ZX8lOQEhSvwZa9g89xqGtKijYMXK1VbnLslcTUDn0d/00mt/+AZ9/k/WjONx
b3sqq0EhBwO17IA//E4IHM8naH0mH5+ouix+mZF2qbJOx2S4QyQml7rfAkeUhD8sjIswd5Rr+kAL
s9qGCOZmPyqJx2E5AjpwPxKPWlqU3aQHk4zwIU2/nZrwWJ+xI94qGPUf00Vy8vJUL42xfX9AzPkd
MQeZDxzuxXPfJUW4jroZpBNoFBfhtfa/t2nQYgQGYHcDlDZ0az+7/69TEJNiA+/tvnofYMFa3wNN
FuPRI2wKEzKegg1gaaxE6BbhuzzPEbU5/5AVsaQGGkJzC0MtjnGNYrIaH7ZQO+85/FrFp1V4eTIq
LupfDvVt5ZCf9SA7lsEGlWoqA/PXsKpcixNi+vbHCAvIX0519AQN+x2Vd6mIii/k8d/EZuAxpD7k
e73bJWg43DWsr8o2yzoL4fsXmlG/OHs29cc0ooJK+cKl6CqCrn9u/oQLz8ZzSUiZaKun4mgDs2Kx
wHEbJEXClkj1ZXJ4GsSS4sAqJwOq4c2EROBATcuvrU8DyQLGEwmrPEQi4fAKCO9uKmV3rAocFwdx
+pSqfjmmgduCHkhJFbtWXJfnv4IZzd04Xo49ubYt7nCch4+OusDAoMMByX1uBtzKpQKjgy3pOcoW
Urz9z7uPc7JAiRk0qQ74x2bfickMOMrmn8JoGMIoQhKABrXOYGZ7lO1qzNY5sm7BAVyLTUs8GORI
/eYOSNI/Crd081RFQOv87ZUHgmH+O+WN+D3/G1ujw9rgjE0r7bZ1mzuk33/ulUbUXooUYCt5jrd8
PB1WACxCiL+a3wA51ph8mIFwp0WLANOy0d+8zvdntZlIY+IPJ8Uf6FQ0XhSVrtX1OEYKXqUfyiy/
8s8kmfNCAvMZ0t5TTJyxa8p9yy99EF7HWJrgPtgE4RZTnJDBPlqh1no5FKyuJAfCI1mXF+FPQ7Qm
PcpegXDdm94whAUzp5hFSF8KOADcq8eqhXzkgUrlipGAtVySOHZ9UkVSgd795ggk8Ccj20kTGJI1
ULW/Ri7E4ETFKJnhmc41jL39j7bQD+egyYx6GQzcjSnnjRrNd3PuUxzyIu/KcKaAMY8NYnnPaqQX
eBgEYLVFcaNOaGLl4UBnZBsFWHavbke85qP55EBsGG84oEMyRKObuJ3eL+1iTDhaxmtliLfTrg0t
Jpz0rxV+G7xRZ2C5bVNf5ctVu/ggodzU4KE2Rw8QQ5Xep3hYIBj1Ujl6mSm67GtooPEd2JRKwAlC
I2N59sJHs+pY3SPsE4AXAuqCeINnkC8Vq18h1gDgnX3R3LZHocQF6Lhyebo7spcJFz93jIA7d08B
iTxyxgb/IWODqV0CwLWRuiOdc30rs7XWPMfJigJZrSvrNHi+21PEC/4iU1ALe7h0nALSj2f0GRQP
+07jGRs7HgbjQvGwj67HxE2aLT97KQKby4Kp0GP5ztE0w0uhQF5xHmEw2xvMRXCfwGjqyLqt1+a/
/6asfBqeFxYZlTjtCCESxbpeQqhAhBdDZyHq+Jm8TUTcp1D5ItLo0JCQnVXV1YudikmmeY4hYu7k
8LEDwIhy8fQKqmHBez5xjTciZb1jaYg4sGRW2AEk/TE5A9BRBK9jVy421gXFf+70d6h2AED4RARR
2Bxqmth3wPbUvTfuCk6Vie/T2/nTeIgAE/lRmMKo79IrV1/iy1px8PPYdQ/6XOKF7O1Ouwkt9s+4
LFd2418kU9Gn/bd8e5V8tBqs/M1pMlwgZCP9I0u/kud+MUjyDRv/Tw+qcHsEiOCqsjYvgivdUdNi
zoBzX3ghmOEk2tj4X5aV9TEIHFj2vp9DZXO1GF8+K1aYeI2egtRfbzn2Xl26vXWhLMxCx06iEgHH
PZF2cnRDH/bNvv8KLEcUhmQ+mtbTSPc2450DlaTud0nDo3R1WER6xnr9L8LaxlZqT6uZYgunLvkT
i5nzMI1yTijnQaMB0EHfKKzHdXr933nwXlp3d5xhTDFTAD8mFREWpx2uk/pQjuDbfPAGB46piIew
FVJiQnpCod6PlJ5xBdfwfEV/XskTqrSvqhGjjJX4kG8SDitKJTYxMcEKfA8oAy72oehDieGMdOy9
MPEKv+VZ0cDzcRMsqdPbB5MvDWJsgb/1SjK1pbWyXv/heCejBEZqJjIqr5qYSBqoFCIXMCgWV+M+
xjFAFn+H0nNtPB5+DtmkBlJyCT98wKUz6XlO3HcPVWChmS9dTUexfsnMbMXtFkhe34rVGZarpOex
B5m1R3yuZ9WbTjwtijuAB1XfQyyelyTjSbLJbWbOukkrey+KyEnhLEoxqG3zuoxvBamvIcfsPcD0
ScoMs413fheHy3jQQ3QXM0ifun0HYvGtPNzWot1hmRHZufryGPqeOAWwPReHzVJOmh+kY5ioQG4Y
fr6VBnH3EpptbnDYKN/AhpgL9tb7GG69wM0RBFU8VxBcsjYjbTrhY8Ls5tHjou78yxxuxL1eoOqJ
HmYAYR2p07pQAem9vfCpCLiC5AC2qBFWEl5Auss0tVdc/MgSrXl500NIbNbXMRhN4FxHu8r8xSn9
9lBhZgvK+EOEtzKypsa9xiOgTfDnJomhZywD3bY5ay5zjiUSqkGgT81/q4qPi5D4kdhp68yAKhT4
rB635V+/3pJFEuQ31gWxNeKJn6JQrvERUg4Ef7pfwaCWBB0ZcE5A1iswD06sW0xHIghNnqMOQqC3
CM/MSplLCazt7YlL0j5c8fGl3mO8I8YyAH1LNCaaQb0M+P14JBYPzCvTfNqkQqHbQ34qGrEUEd5B
GeBKS8nMInkJ9JKSYeHsZrjYPbYkr+K0Mtsj059rH9vNI5ZIJMPclB6kQu437nqpyqnSuJeNav44
uR5FWD7pyPpvNNvaI9T8BSxkVrpHuJWxcbo7lBf3/3aPzoUvBqk+f+YMzie4SKb98z/7BcMCksPA
WlW4LNIKvA6N1cfZi4sk3XkyWI/wwwVZiKBfjOEGtAo9oGJOvfTeIuFWH5UO0e8PNSv9fo095qLj
y1hFjMlqUEYzF3cqToIDgN6psXJpsj/3zJzZAS9hmVzp9qcXSYrvZPQEk0PgbPcOjo5++WJQq83+
Zxm0xjS2s27YBPqymhDx258yhB11wqU1GLqZk9P40kkswNbFZE4ufjSEo3AMMCeaCPb4CpFoCw2S
fxYKUoWIHRmvYh5hvyBwWW9amkfKyJ7DNTLjPjm7+MMdn+FUtj4cBh09C3IK7XlUcXr6wzutiaDf
nTc128jnaMU/ORFgIg5XIU42c1hvmxbPE/CzPyY/pCrqabbnShI7KVO1lKnDJ8Quqqwd5NltJRKe
w7rk3XY+4Fu6gCjMbCYIG/Nv32YbqWo68F8BKe9vEAHXyqGTOO7zdXuu3Kj1HBMsUf01aYHwgk7j
P0Fu65gfitx5ORF/6SYkBibRL4hrzFHTLyjsSeTTIcy8PGdtKfMKpvbujY1oNPjlMGwwm3MabOcA
PR0+SLWIkq1WYkqzlQ0lG0WCnQqNFxz3aeK5Oaz1U6Ub/Rz+4BKOEe01xCgyrW827yTI+R5FPPLy
XCiXN7f0eWCSpKxOzFmgsIW0i7Np7U221MVY+0ykrngYzlpU6apEut577W5Y5V0wfsO1l0BadTgZ
GvFmx2uXmAxLNw5FHGkaykJnuvgE7Iz0jl/aS1CZYL1lkbtbVb6U4Xw/8wO13VT6jTesHy6aA+a5
DbvJ8A8TMR8xYJPP4I2pWel7ajxlLYxnS3YZssUpYprdWaLeBAGRRkEAVoJrbQbOBIP8TCUJnUkP
1OF0C5NHHneXvZz5CsG/VHl//khQdFlVmQFG5NqPEAfdMdHnmLaUYQyaIB5E5D+yLR101hB24ibk
cULzIWDnuB+FTl7MFt7XW7HzUHQduO0slsbtcUtdJZIms2HFSC+pLsdkzqNEbHJC/njSPBLLNUqT
eRSMtFxkp1zL6XwBtihdQFT5se7I4skdXLl8A0+px3+GetVp4M5DWXg9A9ZZ4fmPggvHSNsGAgs8
DTN/K/yUPH8GmJsYK6IwY+tPe3K5hRgLub6unNtRQeABdlvPnvHwWa0aA7teurw/8asIatiEiX4v
WpwZ5XLp4aabnfGNIjEuVzoPS5rvVGl3gEHQ77ZjXReKOx43I2/sXRslLgakGKejj/ze0NaKCVT9
Qqbr/wRd99tiJQ4E/flXf4DDk4LmP+ZkACSMriY+mivgraeN3unRrEgXUvSnorPD7J+4mXpg3J+h
FchmwFJqkTPeVVXbznzzs9Pyze6P2HeheQLcJKNBRKW2Fb/RGqYrm8QYOySKC3kMfxdcchAoz6Cz
+SBcOINViq6x3PDxRF6F0+dpk+FKSXPuG2KtFQ/uPs2uvosz//z68uK0LvDPuhFn7NXt7Qo4a1Ai
y3RXxxfUaKuVjHNdpOUd6Ubp3v9ojzZ3Vpt6dAvKXlFEmAGTjWyCOVhdKMH9I5vu40lsAuXk/qYS
kqI8zTyzVGyl3HQJnTXI02fQU6e6KQY2DwY+tyexoMDRC5TWCPmISw13tsj8Y0bbxa4WDbRy/VUO
zlguPLy4+F3VdGiehNfsKDpvrkUzC1dkADtXk6SDVCDxtJES/nuxp/fwZ8SsYSVCQ3sC8cYmIYWS
EvV9Qw6oxKy1lQwc7mEl65LsHkOzdAzgJVEQTDPUM7Pmk9HUG6lxx/J3NRl0hi8CnoruvKx3qC3i
eDL/F4H48TN56zVdLb3SHeKlbJubfJIx6tMJs14VIfoAcgoX/5OJHb6+PnfcDT7tvyEuZlHPQ3WF
HeLoq9iy9veUzkUKOiLqhqIuuqRb11MGxS5NowfTEcYClO+3uR4P3MU3lpZnNNX2LRlHTMgQw21a
amPRxjDYQea6nXV2brgXbMc3XRm4shxXVCgx1RVM1bwBvpfx39Z5hWWnSuEcMzObf7ROL8k7eLAQ
NLj0H6RdOnlvg2xrLamCD1iuR76XGWa9tEcasNPn7rjzmAmYbAahBXdI6TkF9QalizuGa7/4Rb7+
S0390+aNkVlXfH+kcsyfKq0zq5MOL2+pYUTszZ7HTgMWxWv8wiYIFiSuqsIhhxpSbVmZe2wTYtsz
gSMlY1MZhKBIk2wgbFCFAbZA6kCehe1bdUp3cdLTAF4iCzD3RS9agFidBaHX0cAWakclpgXUgFlT
Bp0dS/C0ytVa2eKgIAkJq4vBwHFbyQIOO0BfI08GIN24fPCOefCW58Bkq6ZqOfXQE+ZtmtP3lnSn
pdqz44/7MRgCfzxEMrtc65uN6NA17aDBY+jWV0tD340sukvBI7h9VJVcDZryeM84kpZ+nxiyhjZp
ZP+dAMS+YuXcPjSAE3XKNvGGL/XZ93GmQtRcGFnZhIC0OkCN/kMVe+Fz4uHWxeaECamjmxYOSwor
88NnEZIUl7XwgHchcsRVtUffv9cSh4OmcHBC35Nv6brglIfb1V3/484vXsL1zdQUmILfOHksFRrT
+MCK+TEkmEV9u3VVyFRpFbMrU95ASi8ie56qGdTBYihAs+9ShskwTzwUa0qbCI4IabDDP7wPialO
KB9d4PU8unC5KO8kSqG0totcDFEeAHF5hmSMnZMu5u+1PXJrKEqSu5AVXx3DpKgPtvWWUr5/8fcI
PEReMaxfNCwRfTa8F4rhN7uJU5f2s7gyLv8WkB8Tww38aJjiIU+og2N2yhi29vgPcCSJ5BX1lF6T
amXhiAbULU88FtcLvwJMK5slMezkbxnw3JUL52SjLPlwuiGf+dCki9veuWwrkcO5WA/kqVX3LsbF
iYhaGSQYogG5CHbuPv4I4PW9blkrJMrQvlXl/ckchKONFpYn1e8gB7awFceHnkdhvf1P5qf+Fzjm
/LKtQ4oEElMqiGwZnD54x4vIWnKG5NHrlmqBMWmExHj9pToRIKJ2OVhEiM/JfhNt1OQ9IV9zMLo4
kvaaam84pnbR4IvylztHL0M/dHq4aJmXRQMiNzp5HILEa8s4hsj5F6VyJLmiRZE6nNipYO0kgEOz
iV+0WT5lc95UxJHPYte69vmnGyJAhBvl/XhFh5S1G1/XdPvkDwZcQmZOAhIw86/2HG6oO9W6bOSD
yU9wPp3hdBZe13u2Tb37Dk7HTx4aOjSIHQLaNpLmb1CpxRU2Qr9DPKM9rFUn88S/wJ9whkxK3GzK
BAM7wO8Z8yNqPDueJ/a+fP6+hA/tiXlDrHj/uoy0aTUUxW5zewZ0gc0kZOUZRRmPbZCSSQbPgdqk
Us7xy949DeFii2fP8DtD1lGg8Qjl+iJfCHaclycLql5cEViD24n6hvr4S2L6qMSx4igCKKAY2uOP
Cave2EvNEcCu3dQ6nvPfQ8HeiTmEIaB+M9ugLbz0U2CCHN0yUaqknty5DJMAb6ogIx68eQMfj89E
vPhGV1v5Gw6AG5i0oBmOKkgaQgyFkCN6eR87/+mXoTy7jgG1RtJ8PLWWdrheeyFhYpshF5AHWS7w
+Au7jgg1FNuqchN1nPJWinKm4a6OVau9pYrGzc9YsM8TPeB1prKYS7gQZlNM3reTcS9xldBBPIfv
EclyONsGCHG2hS1fGwhDkRar4lqBDfLcuqKtY8VgIaB9j8LtIoCVba9N6+38VQqsx4zxpRHJ+myb
RSxd7rGom/19z56jU93jdDQavn+8g/s1N6+9dDQnxmn9lxKHlI+3vIzZxZtILHYh7QWvEzFdQbvX
bULKlSEfBUh7jUljTfVwPBAJ++SleRjmySNvKhGXr6WE5Zf/tHiVshbPc11H7vatbHx9+EfJwjCs
JtP5IMaf7zkHOdpHs0rohEb8Ehz/VvSQqog/BGhh3KKTCeYQwsX5F2zzM1tWclWGLmvFWp8DIg0j
oe61U5E1B2llkjctDtXBranqzfdwNIqqTGHeRtzioeeCwLr1hSVDHX0rdfreSx2rJS62W0kOEOXh
b671qqotRJf9rr1pHU20lGg82FuYxr2PrO9vLi8VnFwf3+stPfhfvDjH+kFw6ez0W5VOaEZTDlla
JY0B9QdFx9Jn5IfJ5Eo5mduRSoast1BwFTV1Eq5kXDU2ufNKVdv4C0mL8Fq/LLy0Z8ZTulcfMC8D
zkh9AymbhhRgSTcZiEP61lWr19l8ktV9juNfAohhnbkyYvNplXrLcLMokb9QTVw37p2P4XnBLMQt
5VLQac6XYQSb7I+DWiuQeCUBQVg3gLRLgas5B7PW689SyJCjhUdFe/nlSB05i6Tx3RTa62lgDPVN
unUlVs0vR6eckdwjbpTP+tIZPIU/xojxarPo/JuumbSs0kZ+GAg9bAJLXoW6gitJx0dFpZ9WhulE
Vgwa0kyZa6/OVgeTKFJpt5a+YCA+mP9fOwIkrf9AYgONSSgX20MwZ0O6IqdAkhm0LyPfADT8BbA6
4e2k6/vXowI9B0K6BtLqftr/yHn7dgpEQg2dST0evQ2e6EXG8pSztD3yPM/neId5KUVtVsV/kuzs
A6gG2ktBeAJEVA2eXquuu3CsaLLl1HKDetuewSYs60Ax/tMa6jgveR+su70E938au3VtLcE1mV+1
6wrU97kim1blgo1k5HW+qG/RrHChkbGI3djzqA3HfQB8pQh9S7LLl7TFM1SpMmTvLPOjj3TPEpfI
Pg/A6qqBMgu3rqWOEWlzhBmGjm1nYyr/98L++bnzM48Ftt4isTKENEPKDkld3Q5jxmcTFnXULg/3
LVNLkqsehAQrHHbw/1M7OtTuYHntpeYnMcQdjuIF/RXLGSQwJNJgJe7CmZcU0ks3ZYCJd6QRpGd0
QH+h8282Qkr5DLiLafbVor6fKgZ/HfJSK1y/zkVUhBfEZu6UkcZn12ss1SjVt6tszzBRDH+90nHu
Yz3C30ikO8kOZ+k+bKrspUo0llO2idbxh6Pm0UkI28KeX4t35pn2E6Ridx42mCZN4S/pn5MoWml4
sM7CqL3yoME8Xi/8h14yiuxbtffwYxmBqzowwTd36EN5N6lSUxZrKLLVUZ/JKLqXQmxCXw9mZd59
7tIvNHFxXPTiK5O2CBiFSc+qEFadA/nRoxwXTOn3owmd7H0sEsqnoi2/A0XzNulz/2ou/Vg0TPXo
j7/dI28WMz10ClomqUjH44wC6zhfBiYtRFiS3hFbOLviGm0Jlh7eLjMiUwYIfesNI6zXBAoVT5CB
is5LaceP2f5PGTZ7CHDfHV9/MEUmg+SfwsL21zko4IlWWcffFFv/drqXqmn/1v0Dr+lNeGIQg7cn
4jzmVeAox4SI7uPoOddSw65y8MOXf0t22ItdThCUKMdf9LWoiphfIc1+yRWTjVXTnsPjVPt4FDKn
77dnbAKLMnjGVJI2czc/ffcytkziUkNPJmAWfkkocSS3VXZgI8IdqWJJUiXnzJskCTgzpNjABSMH
UJgA2/zt824thJYsW8g5+/td4sLfTmC5NgrpKJReCUg54GwCRpWPgVyciNKGArlLNVDeGO3GMGx1
LC6uZ/31KpfosYuwLuTqn8JRf2JrnCbZoRJuDKItxP/kKIR6Y696ewuztpB6JJiFSqhShYelvtTv
BRhaoF9sSH5XLKz/CcvaPnUAB9WeL1ET9uTD7kZWrIukNxIPTygYw90Bl5iW4hmBCbyeEEyqjcgy
kUk+JR15cnmBU5u3uGAYXVDV4J4YbSbsIUsn4eZA3Pszsp84tBqwPrMnxOQe3dHra3kCx00DS0tc
NEWBUcfJ1FqPlzLc2hkNJVIVv1bFM9BhXZ1aJaSbF+j7zFmImD3dn30mOWKzdyHb+/lqYbJcD++f
DXBkHx8j10Ks3wn7V1Ww1PR/sg6TdbdrVf9U4gmb8cvg7ZoAI4GuhCrqil0NVK0R+xBGV2iTLjAC
oWJhGAeMEu6cTABN2xBsxlgEV5HyvZS9XrrrA1Rm0hLqH7Qqhkm0cs9JnPkE3fCJTPhyUKU028e3
uzAdjLDTUp/3ts0HZlCgEkdUxBH/kpV10xLoZiVQGI5YMMtFOvEjvnSe77FzBtpwIU+QkNHr1Lzt
Mwi2yROed2Hyjgu52ZIRzulgrQyX88HR1lQrEifFvP/0LLINSb+zJDmLfsieE9uw+cqs5UBI/rrR
nZXKRnsfUx/eOx1BF2NuHwk0tdmUmZCdHYDKF3lPL5BUy984069eqMkhdRp2Gph+57w/M2UikLZL
FkifTVaphqTGxWCD2VJWERtN79WEyMsCLCOfYpWpGbzhIggNspGiGaF52akFfuVzy7kSyHSIEyLf
lJkvP7ccHN8sEeY7Q4AC5cB9WnB5HexBbRro9n6fDZ98o0MmfUE9ExOL9SLatCIF1FWzdapTBDoc
xz47Hki17CLrX0gn7TyXltooBl9YIm8ovB3XBzeVcfyI9Xe710uiMURtIeR36OIck79Ja6Hd5G4f
x7bX5X8isD+/ctfkbTNhEjg0Ms0br5MqLjh1iCdjtO4UXWGZCstWxAPbu3cgLFktQOiC37+M+Sxm
Rntsxxw/QlpKrMsFoQA4abAVjzg1XNlrYGTFx3FBaP5UmhZeNbLTUnbAKADp4fFOZF0yEFqUhszG
HlaoX0EQNdIxVrPZISS6bAq4nVh3U00h8O4BVglDO6Nqw7YWaRyVq4eCqIfiqhIwmgcp3I3EyOvL
TWZbZiwvrPFTl1A6O8H4PliGQYTnAaufLliB4YHuAE+vLzp2smEI7GJaAJMOh/tKCQlzzqFxITer
P14Rmqe/+MgAKuHtmqzj5OaYmb8cZ7flIif9Yo7AxfsTL3VU8HqLOs9dW6pdXIBh+6Bstoy6gvy5
Ybb3fns3kaSfQJPGlBicd0RmMMQnOm+ONk0g3tVSASyVkAhYDnWUm/6c3muNMbV4ZFDeXoP4khgF
SwGVEQ+AA9NwTsRfHYTBdABGUyc1bV5wdCtnpIfk36WrxuQ8FwDMNVu4S/sUcOtOE7RDa/YbrpXU
iv2WlvpskZnMxUWRUeun6cqnGckL4AByNaDZlzdZy92D47aysXFtnMr6MFp6D730FxFkq3g8GJL3
VZVeUhtYmaXhNDFEzATPmDMwBRIPkSWbfAj8FtaNVOMghjMT03FOOWHkVzpgk7yn78BZ3ET+7a7V
cdJQv/iHBpJBm5Koi3FI8UAf/y4PTMJfIYQZ2ZZtgsj8e/XB+C3e2LqHob2RaS4N87tFiNPXNeb3
XZt2Zpy+Jwe9ful3baiXiX5jJVtHKGPn2x4WWzsRA//bN3glbsdzJ5DPrHwYdbIiYgXtgQAJb1Zt
OT5UFsYXFLU4nSxqqFBrOYJ1bvZrY6Ema2buPktM+pnripESuHJ5cqKyeg58yhjntU8tB5ustTBK
Fer22i0a8kNl3TtgaUHh670A7fLEhXYEiM95NTGaEZ59nh6cXt7mgmMS39FekC0+0duH8mUu0ve8
e+RSMSkBxTsCDpcfLS4VIC3eh4sVmlN4n2i2RLPMV6Sggn9muULmsFydLdZkKHvhrQ3T9jn9qPad
wd06dGrx8Z66XSieFpGw2/97exnms3Di5wEnlt/ZGiKBZYksfa1Y3uw9glwskL6lSryNOzYzKvDd
o6I0Y5r8n+EUWJ5058Oj38bnhJRvwUM+rfskL0c6IsHm3innidBxpqU8eZv/7wkAiw3MGRlKEAcK
Jtn7RFSyTxJsAKLFxrDaGuShgYG+VTfmKJQPa6eC6EqFAzLNIRYyMRG/O17kz2p89Vcz6usMv/dZ
fiyGyWz5ihoC5j6DmVdC4v6VpRqWk32BQChb7ye8o+L8NDW6N5266kcm6a1Hcq3vESmbhrf0tNDV
yKKY9Du1Gr759UcpY1j0av5Ot4QRVRy7/vE3o8GK9GR1sUmOynFvntJXWPVpQe76NSQDftZQkHjJ
I5vGTszUYu+wjw/VYYV484GCvw36QGEN6nBI72yRil0gkRDDFjnvtiu6NMGWOhAKs/ZzsJ3XMxkw
0iXCJlA/hAneeKy/ZE8KSN2cBF8dZ43K/zsjKE+VtgssH4dljKYqyxwEvWk/Jy4DsefTSBXWsp7e
0hGWyZ5oO0j+O+TolwZV8wfLQnmh70XCllECUzElsb0RO8lSby6OqxU357VdhxRAwbTyO+GgDaZN
MSeZkcjB9wWdErTX8KRHBPdJTy+BaMAJooojDNAu+ObVZKRwVaJsswy9wmXgLUIwm3b+mpvRnJNA
SV3rOpgFnklnbkikl5lxGVLoAEsKoCmXGr54d7KoFv+PLX/RszNANGrgXnz3HtU+xAll4lhbp/49
TCJIaNXsBebjoJkYPsrKz3841fXo/E09Mt2mBiPS0s4+NZRQx4WkT/PydzSYzbTfMy6wVrkxqdRC
OJTCipzpYeOK6NXP6luJ+txQEsWoSmbBXQ2L5gXm8YNCDMuS4GckHrYQcRAmXUI1iCx4Z7fMY8lr
VSf4rs3V1wmh2f/4xE7jbhnx5bDoeZlx2bqvGvBhhY9DS88fFZ7r3gbUUWAWyyjEKqnhGNJ7TwJq
ZWtdnFsYK/QpiUf/yrTU/a3JNItIdA/Gk8R+cxqKImyJxzXe+zcdA5kpD5ICAhS1+q5MxdHes9UP
8CJjNmoqb4J4INvfbS3BU8BKcx/sNySttgss7kNLBkdTH4rIR8Eybbvjzo+qYsHIR9v9Z2DYoafR
fzzRZBXXx65BiWkPXph1x5KlQpsRYgfyweGth0QCfFZ6Dk8yRB7qyGw3plyKUqXTjDn8JBvHlgnj
fyuz/5wCl0tKA/Qxfu3pCO1eVy3aFqJkcwze3McggNbsttAgqLcTLtgQ9cIxpQEMi1/DsCvq0MvT
Zti+Fymuh7LUPF7upH0sR8SDG06Nz5pXYVBVBMMdLvJaNqlXeoPsI6McKvEWdg+/dE75ceIzUiiB
oKZk5s9reeCT0Qsb5U50bWEmg/aG22uLm5vAg5QMbt0N8ANF1raxYeM7qwgZu1FsduzxzAAyKd47
L/fQsnJ0dWZ99PrlP7iLt+CV0afYrfPu+ZTqaOBvxpU7Rcy0H7h8S7Y0jGyvqDNE+jK/K5uTtYed
FcUv6McxJMtAyuhSFBFv3tpJJw+TOXsBtZ+oQJ7WO1XTiHJzAu5au+tDeKOR6N8mRAToeOuUZFiK
5nzbbb1ynnwepMUYDSnNuXXcrf+6b+of7bgI6Hm7hVmickqVon2EoDAhaPGB9wY8U8vpOe/VRHdu
K5O2eewZK9ts4gCtEnHFwOB6btFz4oanrV6Om+aZ0hbawSVJLETdkKKdQvUFgyEbjeSe1p+ct9Gb
4dMOJtCAT7d4eBj8JmavT5q+/j7gxEojq7LNufvhLZfcBdoIVwjt3Kv3FVERXACuijdcd/sKyYOU
Fux3gfN6bu4xpb8HXdJVFkM6EkaztIswQMX9/76laNxllHaUWv6iK1O73XzVvfXT+H4Wy0lvknoK
dnZmiIJbkRPKZ3rVSzP+6iTzjxEnbV6U+c16wkhsTQUrxwQ+qr3rGbGeCR9mA1F4U3QZek6FlVGk
jGJpA71Sxo8cLs4uHFJfqjzSvC9fdtRkFWQWVnPlrCz8sosPrC0ONQk+C3UVgYKkdqkAB7+7EnIF
8Dn3t1c1GRjOMZtHXCsVjp0JmTNWd2RFynnGhSEh8cEruCfPF2DGl5vFUiXpyWRmqLgdR25ur84C
3COoHd+GGtTdm8zDniazI4UOg8ajoizxQ1Q1JnMWUP+t33nsHANvdfbGDv7+q7VjMyb8PgE9QY9Q
kp5F2/o08UppmdDyYUqndxvNhYtXjcB1WxpWRc8ncJarV70bNfPE/JIEi3e7WYHXj2R0cof4y5Hj
ZVOvkwt5FTaksrajAXX52Cf1xo6xY8Yx/l0Pl7/AF4NJnAXSIYYhP4tESj8xkJ+dfcvGrS+766UR
MVwuAdRQeOAsqPO9UtkuUmA59Dkg2NWyOJ8SLbi7e96bBN81UDOYhfEvz2Qr1k/FjyL+7smA0cdt
5IVZu1P+38j7i/H+pC+1kpaxpo4/Ii24nwWpcRj/lK9kjXVqAuvXuBP74j7kk/C752gPB/yy3Hu1
M1tvhYfA/SH5d0318e6sYjfAfk5Ps86OwlbJ2zMlQl3Jqp+wKZ3serYbI2pPEMbwQ1FrEPEwaY+r
i+MGMnEk1102NlflUE16YOAt7utaXTudPba561FDI5nUjuax6Bp4ybLZplRn5KanoIkOq9INtyAX
1cFTJNyHp1o6gZqsTZojVOkif5OiPwmiUB0NYS9zxNJmpY/O4vWHO1Gttpe0wTeP8+CZlUjfRex/
L4Q09hqdjKEvyuWNasK9OMb5y7ETw5T2yG8KOhuzZjVX8+eE+WP2pwnccY9IhkSM64pCI7EIEQ2+
UtLa51I/Qv2+MJO5IZ7JfqmompVfmJLzqmrrXVre3V9POAbQBwrdiguZ5pUS58dIpuyL/hq+A1AM
ROUmjQbUhnyytlklQZBsHlC47X0LZIRGwHKXn+Xj/m+oJ7Y5OI91eKsoJXwWfRjwaix7nnvpwSU6
uPavwfakD8YCHgFmGAHdzRNZTmxZ4Sn9yf8QadgDxAD5QVldwYTmlZ/qhhDYkfQ2jb2jvi03VCpM
WufFOE9QVszaX9CRw3cWaldmPlW1i3LyNGdblNOW6zjS/gPa6TkKDEaCwY+O4Ub1LbEKQDedeSAB
7UW5wHRi8x6kZ1uvY7CyH5uBhbFoXO3c5MD7BcR5AXrLDCYYcwGsMaKrNicDfUhRAqe2Srijk6YG
DADWO8za1F3Qjn8utYcfLR2XUoErzF6Iyy/5MafmcCdFpLbr6aNKWOoBRq0Qi/UaJXWc5Buw2QsC
UdZyoz2BuiVSZpOzBjLZMRhi4fMhGlIGokoGJS9ltGEpHz826fzHt3Mtg2NMeBR163kvLHUoBA7I
SvpUklLz5jyGBtq9G8HnUsQM+W0gtCiIM9E2WvvoUmEiJkTeNOtNh6aYv91OM37yUDYGnyHk/BU/
1mD4iWTDoxF7hQtAMUhcEDsMuEXwYaTVsdHkrgmmzCavavvjhWFpgzr80qSsTs1eL1D8QXVAhoTO
060lGh9pRgFyzSvs3EOgCE18tZFugRYhyOPL2g+k6L8c+vVVMTQf4jPhH15qEmS51TboPbIoHfi/
ar9RSVD7zRj3xzFcFlQLVHOVIctjj5kf2ik3eS/+TOFmYFNwqogudFPxBZfUpS+goclrzrhSlpQ6
OfiaFaOEdqHRcNlgyA30nxBxo9OKTac/KU5FRH8S2jtwWKyk2ZSipHI6TyQds+qYQ6pVuPAMYPdc
4r1J3kPSELHhfi3pcn5VWpvWE54M19uAWicfY/eCVQeJpIF6MqTn56fKVXLOQ0pK5+evFgmVO5kL
XpqhrSnaDGaH78dvKJ/RWoaRwQ/k9FPwWGWvfKTdR9yyq/hsim4y6DW7eu/WsC3jEyv0Lcw5QjR7
w6bfOdV0M8XwH2rqev4xR2Xgpszdvxh9xRT8LU7j0q6EaSEm3Um7Ohn6ZI0ZNLE9jU7YfPjimv9S
8tdMrGp6hI2wXpaJVA8ji5o37HjMbXGNO35vkcCoRJUQ59LnI6J8qbo8dGRuy+AfbQF0KW0u8tlA
D4mNQSaMsInN9p37hwV5XirD5yTZxmhvKgGO5RhCuiUderA9SaN6YOdXms/Maake8VXfB8OzHDaS
qxNC4ZYf5vJAB/7YuCA5JAVeSyLy3fHTBxdmIoBKQ4cqyO38JNV+7YvloNoA01G+eOkhdBj1qT0S
3UHxAbZ1jLqL9SQau8zhZE6hmC4aIcR18r+P40bG6omDiVvQ8vFFUGzNDpwHIymLblltR1j1h9nC
Anc9zBvO7FceKJl6W2kAOxW6WsnJ81QE3ULVFTN5svuw9tpsroHgBBP6mWH5ZHU53kuuuLuXocBW
6lejLWnE6GkPKt7rVVYEWgPukpr1fF2WQ+t13PwCWZeQSdFQeGDCkrXvl2YDJj3YjbLvQegKYTcD
NkMHinp6lpQSBRrDdOyfcUoskgV8hda44uGUigZ4oIoNMLIeb7JD0MgcOefzyqUWa8BzSSd3OGnn
opxY3D93wU6+WQ+MpE+bzL4gae3xy0acmJjWsC51IOCIjCe2goj27M3BOeZltXVmKvGOkF2olLH9
z+KwmBoz2CrHZpYw2T5cwCQfB3J0K3xbi5dC0ZhtvEhZFVTKAnR5d7V6rfXpqegUp+RVzIhGwGXN
WdhbrmeXB3K2wga/8IagAIBIyld1HkcVt3gIWEEFtgMarU3wItbt1e61pyxMPPC3Smp2rN3b3P5J
yylOSRycxVtYzqXN2G4TGulw1EWHBCYCxrMe3KvfizeMwpkslTmYKE5BpjuUcTU5/adkYgDL0/He
4PrXbUNHacgUk1IOWPecB6DLO+JP2IWjE/4qMcORSvF5jVzvixZypy4T1f+bWoAxRSWIcLVOvOpc
JEPhPUvwOOKyi/7gFHPgZusxeCMTZXl5oUOndx1L1R6QhVpTi+/SXhpQqU1+RusThi+kFUcxvKud
xeWTycELBtJxLy7Ibs/oulIAxcAZH8RNnDkt6l0S4LCA3YV+MAEBe9qTB0ipOJzBuo9oxcovTJnO
u0Kw39YwmUIz4NxIa36wiOw4IfLUkQdxaHLoIrdTKeVac8Kylkv3iw9sDBn8SS2MiJoh0T4+ZlgM
KMwO8NdSBZ5q3z3nbXg5R3Uw/BLJ8NpMNifcEn8fTUzU87yoRBsqKMd6W7lZ94XT2lEUmRtiWB2h
gUVcfUWk8sEKxPvezpFQe2lhbewd2T7igiOHYGTqHzAAzTp/fUvPLGZvqTpKCyNkxJEyiFwcDVTJ
whQlkAZ0RQ6NcAtvn5RIt4P5hF6UimMgaMIgtsuc197Z19b5di0P/aojJvYjbomrJzsr61wyDukT
RCeBxKq5XUdI7IQhwKbatswTTzEPj4YpFxrSvOBlZzCtLwwUOKcOyo2IVNaIKvX49rJcJvISM3Y+
gtVWXR4em5XOomEiqJcagLLJPTfDTUgqIxxFXkuVgrcNsol3Vq2CmQSYU1yu2Wpx0eE4tGJ3/knO
rgwLPT3IBmYEPNMzI6ikxgXuQ+MtgNyPt/IMQbBL3RRaG3ZakM0vfUgFoCH9l1/iury8Kk28DgiE
PEyySGn2IePdfttMl5vH2cnarmN3npLuN6sdgYdYaHI43Gg/s3FY6B2ddZddF0ncF4Hf9KX9x2w6
5w+f/z/gyjsyzOzUXgi6EggXn1GJPRpwzPhLq3C17KRTJLYhaAxjGfdZbD8iMsVjb5ukGyurWK6v
XZ0SzC6h3zN2ZoRuXm3SCMkiXNpmxfy54xOWbnkDMttfP8h3600M3227fjkzLsPTKhIP2rE641kL
NVpAvKEHUpNzLIvrA8E+hSWcn51+Y7SeAvs8768ErsSf2qqRfmUPTEhTBi6ew8VS7qXq+EG1AcPN
HK8DdhBMPmlwqpAWY7W6evuQywd7HgKNTUGTT/S+rRRORbTvbcA8oJ7+p/7WTugt/6jTv++Giup5
wcK+RXFITshs7IlWR8uRbAs5b0AZyBgD6nsNX53ONoIjFSk3a7VmeHrObeaAZHDyrwRw9dyKjCIe
kPZFghSromPPZVTB8XJbBzeV0rVuCOmtoTisMxdqIdOiewCNnD0DYlqsNRRMx44ue312WlLicUOE
AfpleOioOg6LQ7AUomXRrisxwKm1UUXPCGzr0DHSefuJQ/1JTl7eWsjorPxVogGn3bCc3OD7T2NU
A2IdkmbVEGYcXoesfs5nJT4K3+BId31Z8dtQdYqW637FGzVchdR6HkIirlIyQ01D6j9xH5JE4mn9
/++BLKD5oBUBumuMD65yjoJaEXONtJI6mAvnDbRpkoqnBQEe0JCTUdmK+zl00+995nqVeqPBOC27
Ttp5DjdfR0oWQTyfTkY+kJkbkVrtrMQ0S7s+yyeTmYWRIC4aWRJ4ZIq0khiVj/6YdIqBOfSd9f5X
ZdiAsS7//uwVH+uyoM0uBAP+pbw4kQEUxrKbhj/eIioVSBEJk4kX2qC0qZ0LlbvWmGQJGnueDlWY
VhbhnmMzUjRSbJS5WzB8UH54fzNIwPGPg2eFcnApPk97nxxUhpz2BJaHGpsMpxEi7w+C+f+vpW/8
ceeWejWs3G+bGSnaxwp8LbhLb36t4lqlSOlgZ5e/9Cd94b4j2R6KEbqIU7PUKlB73mlr2P9B/yIh
w4WBzFSXmEXcSLQESsxfJnb/MB1cj+IuAtlfC2IoZvsvDTjgkhdbDkjNaNYsmJrLb6z5E3TepNF4
4JbywJ1AnP5S2msBQe8gfpZnsVTRPln+ubVCjJcam5L1LnhVLotIge3MZ3ft2UvhW0qe/wfeU5sl
ugVdvVlgZVL3W7Cm4shluTrr7b3d83VfFxAkLPhIDoXheD8rR+OyFv36Z1j9j4NpdhpzpT+nz02D
BqnkGHlTCqJ2U5r2jYj7a9p/Jf+o6JQKpjJUKt9hu3pj47GMVK3dj5BOkl8VrCgcVXjiX76RHwII
HLR3gjZ1Qn/t3TaMbBVP4a62en7CYVG65SvgG7/cVaidlH7AME11fKtIKClfxBxXAoU85ZrKrniP
4jo++S01oZfGOwZqKZjTK7/98XVcUKxYnDYBTQ4yKeWHBgiHHqCwrUYB91UGceAThJg0M1evW45+
q4KQZIP4kyjZcMBpnqPrv7JEsPo1apV+C91rIyUAXrRQxBgog7Sh2bC/pFKlwzO7AQjTRkqyYsct
GP5h2hA3eMVuqtNvIVNNtjJl9Hsaebgku/ftYy65pmYSSpow2JHmzFI11lurMQRSViRWQMNKf/uN
rsBQEW+scIIkWPpl+3CbseLdqrDWxwTVYlsF7bjneA2Qaurm80N3c8AgvHsY88J8MYeSwjJ3wHnF
4FmWb8een1s/kTzxTzJ2jAsHlivx/TTCKZ/f9SemZDV805VD6HSVBKIhMpE3uNwTsK/dX9lAU07/
1b6WMbsc8/w6SA6jigkRK7yb/8J/xFQQPB5JIxUZJdMN7R6K51jTaMvyEXEI51eodTVbceWGifNZ
iBn/R0Jeq17nKFqF69U4u2q6vCUCjS6Q5SLsLOEyWyBaH7TxRFCWtryeZ8nz6qBKnI5uD4gZWvSw
+6H8XIbO79JC007ppG8uJd1YyV6Wp13q3leMYF1ol8KjoAxGRKqegeTzDqZfTTbgg/jXF36EuS0f
nsl+heTwI8nwYw1h1S0/IgveNJnb7X3fFIBO5MePeE28NK3tglm/C1GZCf+z0aYruFVgEoNbp1VJ
KU/LLog87YIkQJmbTdIpyaN7hE1lFI2/jmyu6EBRyAz5p4BBNsAUUGZovFZERUkl3WGv42I8h/EG
lVGVm6QyO5S0Xx4TWZYOw/Qhj/D4+nKd7/AviWWHqlXamfHjmud16vBpqLXqzPSlO7YGdZEfbk7w
2mSfcBMYhNMFgohzwbNeqfwEbrJdFyXMvEu6iQnGhv0/npoDmIHPdzquym1sXk7iXoDds3Ca/QJP
xB+y7drCvn9EFDBezS5rZAz1fdRcTypc6bd8D9BDGceBIURfmjv8w68QOeRahILuv2VwDdF7sXj2
e3aMmsY6yyvtFEtljCVEiCRjKItlzQ8cmYs6RfLfSf3O2hXRL+Szw/e2wjXmhrK32dBPZzG6ZgjV
qfWyeTL2hui2px/3sTayBcuUa+PKYcXDwLXQIijX2HKJrz1jiqMbjipj9F11kf9y69AOl3K/tYjs
7urCb/iDrWu3WrwfXz2H8c885oL50f5Um/7RWI7KOJjPZBQbvTXi5+8xpLhPdBqkp3B+zq6ak9nx
Z+r73yruMTUrxoFspB5F8zQ2wid1zjYANyhytLINP9ErcZSCBhBNs0Oihca1WDkUj3RGlsqqeoc4
pVhRHKjVEkWEOtJyqQFHCfki5U2Hsulk/CDQdvo8WPw9ea9Pu/lYBy3VW04giQZyGoyyKypfZzJr
8OQI6uHASqNKJre0CF/S2d5MkggpvnMgwp4zqWdRGuE6Nj/pCfvxcTX2Nd8CkUvRwfrOAIgrxx+e
FT4s5LewrtBUx2+Y+NZrz7Wagv3TfvL8vyxMjjYkv8ERfAwWvDLAYvfVXVRoD+hxCNdKg4BIHoec
hfC9036LDxXMhDqIfJUPcE6dOEM9qIqUb3nX5sPEL6JQLRJtE7Y4Sbw34GRXMGFiD47Mn9lzXs9n
z7nPxfkp40HJ8R+Gk8YS/Els+oqfiA1uKO2e42g97ppPlkOTctOsfxIy5ueZVNTJZnEwtKfViLQV
I7Am/Qd5YSW3g1J3WG1knuBpkPjX3BadLRn1ajPyvYNbZFzUZq8QUXFb+EvV8QNk/Ox1kmcKksdI
fniGl2RgYmz14FpIcfAELd9t9h73ZpWLpyC34RTX2lFqP+/n11ydLJ0cjOzYX50TUCDR0ngJu8/M
c1GzwpWN/wQnSNPqTMX+HaVfhc6RjSj/LK2V8DEBGRoPKhrNCdcp767M0xQsp8P64cZxz90fP2XS
kw5l5bCMAIffkuZpQWMzwmUokwYk1ph07arzrYpdeTnRW8VBfwzrPI13453Ez/XJBwCfzaO3BILB
x2zm4oQ0i3A+rZD+/NoOdLfUycJMDvzQzVIqnEpvEMn8iat/s4tcHvwBcwQO+0ismc2DoMJ4XW9D
5cxawgGyEmTThI7XiAAa9UlOsVRRrheMRxWn3RtVRwRW/frtC+KwT4tHno6w+dJKmRg4quqt6nfd
zJ7tsAoNq1HDMGxk3fpXZB9AlExxfeyCyBg6nHEl1NMtJO7B+kyQERbcHwH47r3q1+KUKPDnsz4K
S/9qZR+aoFEqF9ILupMH8itDwTxBTq27hmmyl4G2T1KZ5gZz/jFmiCsJWkRTNGSzh5H+278OGh5e
LsMVaTi+qqgnDskhobqpxR2BbbkfgyPI1nPSxKv63LbhPeBkNC4I11CCOLm1cgiuR9LmOAwCnI00
YMZAP59PBynr9E2nYKxg/uQ0gm9LwJ1zieHGGnIDEvLN025AnzOGjMtg08G4N3ov8RolDqiBtq4U
MpfS/9GBagFthu1+2T72dSCFP0H6JYxJgUw6OhQnizCiFyIqODK7Y52oUPyZY2gX4BqGYA0kzrJr
eTyUgZjkJ6y1PZZFJmLR3zZq6xO8lOPhDlqMufpyuVuHyPGr49Z6tgd7Tu5pFG+4s4kssdzIi020
EY4kq6sxNa2HVzv0Nl9HNrtwn59EHs0Bq1z1oGPvGLKrc0KREHe3GffMJex7tvM9AHky/Y1rQBfh
LFmDkENduHGf3pZGGwdrYIVxRTjm3BBfjlOeN37BfNnbEqfRDh173FkgqIrntsLjLL7CurkcCeg6
/qIBDL1T2b5NY8kd27tb/zY2c2K4RkX5DwI/56LHBtY0w/N1lyUmK/8Gwwy6tWuyKXlMWzlDnwVd
ezLuBMIjgjM0lyG4uPcXgDbRw8PYiJRCuk6QwxYLybUhG0z2O/rn6JwD/aK7s4XQwhGBobakb4ZP
VEP4PVQ0+E9KReql2wxYWodzKp9x58Xs/oRDnlxPAUxHErTLqohxf/uv4ruL+i4mPp3YNsYgfzl6
Uf5MC0H4OvlCot16ZsOCQ4wR5biVHXyk2/qi5S3hSPyx0Oa0C/+xX4R//BiG73LkjVLBhufxHC76
ceE3eKp/s0Mu5SjOkQ4DA1JOOqTIZ/9XEx3C0TA8XdVtzCDCnQePR4E/ifMm3SgcGGto1nVMW9g/
GvFgXoXjS+6Fgz6mZO/uNMJiQuh+jzWLesnhZt0qTiL2tZWdCGdTog+m+1yEQZOlwR5oBEfrICze
NPpJ1TkakSXp6ZGo+JSU6fbmxxBa5+Jyvu5pF734rxwmcR/6aSUT+mC2SbJuMppV4+R0Orc7cX8I
aYmhCk5ZFu7FXU8xzlQ+JkMbdy+ImWKFfPcX1fVrTYUvoX4HAajWhq8Kpd9hgVqD5lLe8jICAqRf
P9PlUUyMKu2HhjjxMhRNEx4751//81Cf6aG8zyHPI1M13vlledvXJvVpYuHCdZ0VcThmrT1HRLL0
hSr8Y7SnkSTauKdyGZdetJlDbtdQwDRUNU3bYCSeL8nBYAAq/J621UuXqysUPDodXjxhhLXyZzQV
8NT1gJvBS7hk1hr9XMTTwo6BKYAFDyxftXhKAS9cYJgFR1DbHqhmY8pzVGylFR+Ildpr6SIl0rSE
SuxDH3fGE4NLDOcSfb2Bo/9XCp8ryPe4x/AOWIyPNEwffha4/blfP55g3a9dy6hBcQnSjopvAWs/
e0Jy+sbH9Bm8uECVSm4iB4eggD7vMvbIulgAmpTCdvYIp7AGuJNTojhsUsvwqIiA5w1kiEF4Nke+
8ptP/uiFI6KAP/zUKA0dUllI67sB1Ezz+oJEnbbOlDlJER1tSiKg5YZqIlpUYuTgXRQV5VHGvG2W
ao7uTRAdWP1OhO1zSN5f0ld86P1H0Q3q6h8qOl+cA7hkcGrF6txqBLhBflMqzFuC+k0pEog6waZ+
xn+gwpNmmCi8ekdhdRwq41S7RfI+aT2OOQx2QzjrpX6MmeX1Ey+7dFYLs5qrl64y85f3glChJd+l
ta6fhqf/vDBenTn6Gf0npTsqFY2559n8rOCcXP3MCxrBjjuqHxt5/tnaYmnI7JA2p9udtbdr05JT
+nQ41gakLq9Gjrz1fWklu78OYJ5U/6puiP1bMx1c/GyBipiBySkChTg+xIeQzaPT9lFGOtGdYA+p
c3WmNhjN5jrT4hSVMZUDeIIYSOBYvw5XFD/XB/CRAVLv9LIICjMe5uTdKg8nYkANTass4cnKlFJP
upaUigO4QIzFCXoiQsh0nLY7YtDxr2dmennWlBqreqSadwh5Dpnz1p46vdk5/jZUjN/LNQLF1wQU
G01KA9+lDj+qItZQy65zDdGxBtciX3qXSfir5YFP1zmxvgw69AGAUPtze7nzwp5bc+x+dz/04fhh
PiNk5BIqgiVLPy/tXfPGld9jYERMgFIOJxRJ60TqUAaD2FneFLiEDroYsOWrOnEuJRL2hNbprXcg
O9wkJxb/w+fXUr5hNvi8puqTsFqQQNGU62RQ2zGaf9MXejjep1HPeEfg7bm42urDu/o4j2Zua1FK
Qss/e4jmXBsPwM1mEQkbUgcKafLyRoBYAG6p17iXmpo//9PI6UQ8s8McqEr3tKS00yLJHW4fddh2
gJYg2+F8OxqhXWCtbngGyq4IYg7b+omYrXayddJPce4ApOYNpAEcSExg+1x2O6TrAeaGBtJ+uf4h
QLLIjRR3QZ9L1/CVY7VwIcz4RWnthU+5kraOUivEsxd9OszFA8jmXz8hVlUw4/Yu57owqYHEaHK5
vgNmmM+K37PuqNd3WMa4UoF2/8XdtpaF9Lil+etldp8SyGGNxlwh7xjFHCR4zsjMIGft9cMCbxHX
r1X+ztbfPTOG/D76M/WaF4ecLBlyfaugrMVfX1aAXOnNsvAAVHzqPdM4MbszercDUhEhNa69jUjC
frUgHCFtfx7Pzhu39AVjDB2wdySH0QFvyurWCRseax6XtMcUpgvxvRf1VBwWqFm4NSex57L33k7Z
Ss3VF5GmzQq0PFgZcStU2IV1uOqNz1E6Q5QFVbXIrwzsNGuQ/q6ffFa/bVTJt7bl8yPM7NJHrUaS
ni2zil3+Ep2FqkTrLboALJ4ADeS6akGvBEw15OLL/ZCkZffu4r64lggbKoMl7WuItWEkpUwNW1IA
ZGxm8/yGXjq8onzGKnfgrtaQk/RWQE4sWKQ0zWuyovwGmWBoO+2TSS8F/4FYY8x95pQy7O/sA5JX
VBRV9/P0W1xxZdj9WzROcIbkNMNEOOvyeJd5wBa/qNlcUOApI+mcUjla1Q/sokWkOBVF969sAU2B
D0GnIj5S1Xo8GokVK33yAlFMIIrbRAC6gZxTEKNeY/nB+m6tnGPU55v/8tkreO6kWRHfUjQ8hS98
O1u5Si19I2uJEA+kYlRP6dV4uxgpS5wf6vWUzt+9cIHfbkj8U9lNi+t3TgyyK6BY32s0XtecIluQ
Hvfhi59zlKNaDJSIngNylf1nOouJ/A3SY0IDX0PmFW4FQVL9Kvawyt8wZEvxV9RhujBEWX2JOM4A
HPffjary6Ro44bN7ruCtoMaOqpKdL1tvDfxGArAY9YaybdI3EPq+jb4l3r8heMBKm9wZzI1d4PI7
X3VdNDf9yU/nL6L1vs/mcGgj03BGJkUE0eu6o2ADyao5y59zYRcaXeeiownxzxFHdrOv8EXDBUzR
FEz4YlWI9bcCu5CbnD+2Q6NQWTB+deqdwf1kH64/yku+bH7O+uz7Db+43Qcoe4rBUxiV+DL8Lpyi
TqcqwiGaXDStr4anWUEEVzlR5Isw5j2P1hQWEPHASqmcXfuY6jCXHdbea+gBLUaHybCn/Wz/s/as
R2RA4Rf8XNCLRanWzORPWN/kwY0N75Kkif316nhBopCB5FeLtQIfyTMGmyDZ/muEbLQpXC7Iokdt
NECjUVVfvUZVYFPD7dH+1/8J5W9AwQBcklkVqMFVthp8vA4LprUJZb5hRdDBHQQBoUA9NnTk7nZ8
XAKkDG7SUZJgNu/1UVIP2YouHU8jcjhvu33OL2kNSMZq/seCyjdw11fJdzuSwnKX/Sh6tSVbr1AF
MlWU4XnAByN4wKWO+mUXXq0V7IjbBmBgtQ8pdjvGb/QbmD7kuel3jrla1IeCmCNiijzphVI9paBE
ADG9AouR7nk+5zXQXiXcz+TI20sf4s+z005h3WEqDjWgKRdmsAn9MTLExdNEXkABZ5HfjFd2c1ds
M0UoEx8Rmq0PhbaZpDpjRS69ORKtJfF66fcP/QlUi7Cb8fXp46WvNy0JoihLW9deeb795REGm8q1
6sdH+Iq7YC9yGxtdTt8veKiccd3aHxO0n46FE3eQUFPl433nps2dqwmOZfNu/9ylOyYlg7YCKu75
o0GDrqe8bV9/DU/fyVLdcngYgUpQ+Mq1T0WVHpP6cTTfRnpYJL8PGwLEQvN1XEcd0M9Fwb9fwZVS
7vrzTrXWjTK2pQEKEy3tgy2O3KMLVuywmPvWR3bsOK5aJfAKSJWjgvvmAtQumusLXrXT50+HaLO3
JFYg7IQkrptjgbwRnouCS1BOeIyESo9dessVNuHTdjGJ/m/lsLnh77eem3/r7Ws8MQFEAHP870n9
148yNgyUAzSr+caPRXansbHj+vK9e2nEfzyPOsEo/p7n+02ALJEj7CWqFzV7wqDrO1R8xpFNEmtY
r54LD8et6tRK7gca7itggTq0C5OiGhWT3IThLAZgH0D6q492zhRnYW7GIsTHPD59mw9claK4TQEJ
gCjZ26wQ76fH2IuNwF/mRcX7lvGcJoSyeeC9RQ/QCjrm7cQFW9CuBzyIsqsC1I4nAy0nYRiiiR/I
TfIXOAyV4aMuAzDJ9o9vJd48oa3Q2Lp7iwdhlkQ6iohYKe3HbC1kFtKxKVa9uszHJwiQr0hfFiRj
4gb9vnwRefi25KwSLAoo5vPHJLkD7fzyBBzUtMjORCOgFriJKHcxYclSHqJ7ncieNFWJyPHMQYWi
pzj7uQYI3sto6Q9oM1AhVCvHzRny/Lu/Sjt2Ufv6v696MkhBefWJ0uRTjKz7/D2NxVvPzyH6ZuJ7
Dge5j9RvXlavtMaQYcDKJctduClwan70OPXQyJRqDxhEFPiqOo6GqmxibbPOHFhYBK/YL6hkfW+x
0a8bp2kB+j0CFCzrqGh2D7PDbwX/gw9SLYpDliJVATe7HmYpFk1ufiVC8hNDxippMhzjb5dK1Com
zJ3C/dgGVkI73gCXw1uHxif8zvIbyZRe6EGR4ddGMQv//iM4Lg3Ufxn2AOmYUj/WMGwzsDkkigLl
vx8hSq/xh/bYw+zbbKHBwxlkxjMHE8Dvy3h7FZPhNdFe8PYQIX3gHf4dgUgN+uiVn18XjZ6zJTHs
MUsZ6y4ZNZYVpfahAmby//eBVSQDp3Zm/jXv8jpjMg3ntLiODBHnC7IsewOAm+7tswSq1wP749pu
4enG83b0lUu6Jbz8repS+T3deSMH2WhCSocwcs2p+S05V7gtvzVQcj65QayCf/feH5317NX7cVg3
oXohnzVWc9de7xxlQwSpGdI8mT8e/olL4lvzxBWWQn0kBPBvSn65lRd6Av4fPeY8Dfx51IeIkD2H
ADNoNnedkmxpTtIfsGAhHX8fpCsSrWCQ5Uk61vZSGXQt7giDyrAO3LRYYYgYMmkRbFj2ZLdHud50
J2nu2H7nPFsPYB5wmn5b0vcpKqQ5XlneJgjDneEBqkl0wbxzjngu59UsgV+VLcjCbY2kIqMQ66ER
4qYP46Zt8hkuQS73cb4chUG6AwzrouF8x8MJrF6L99yfR00Cl53CNgxr98s5ANQrd8eI/PjRaA3B
6a+dA46T+1B2+oh8QcarQBu66gicAtU79PifFqjpq/P/xmuvUSPyY26rBaftNwEEa/o+xGuEozVM
h53jV0fhc4CZhZ+xn6AwxUqF+nrTPhMREDL0iOKEE1zifRTvmoYTFDbKN9B/fKMCVW/RwhM0e2sf
dI7/exr1KiVdhvlL5ogpwajZTJatPSWn0pRS6zkiYCSl5sAFEJAFN0RLmRJ7QucAf7ywq6Ilb7a2
nn0mEePq90bHXL27DUbWoe8EKMUP6hwD2LeuAlVhGOoN5f/CLZnP66vYE17Yk6nK3qlBxUYtXtkw
R3DLWxFoPJg4zQkghzmAjnLZmBuzqPZrJjxLDeDyj4q6kaDF+UQgH70DoeZoMIRCg6Ln9ZPu6FnA
+SiDeKPXH5/vDVBfTQ+f91/a32hbMudxf75HIbLuI2CYIxvnwlsNWke9ipIfzO5RpkcVcE13TLyj
p6ZCVCutdQaxwfpraAEsJ6yw9CzBqOUOAVMJ/AMzbKlxctzeH7cfVaK561i0PDao/U8OIUJzbLOt
gbY/I9vr6+ldIhnVk8tHfOb0FY7G+3xmmQsHNnOWhJlZGxUGUuBFd1gRhJUR65of1yFAuUq6vGDa
h43y7uKA2OQd7cb/gsktP3CPNV1FQOs2m40+NSqmg452WNnO7LoJkGtfhhRAYMe8EHAXRpxQAjcq
UX0kFu5FT2ou91SlOHXt9VOjk+lI/xZ+Z7vHfenSV0Xp6B0c6zsKnqv1yr/BYbquAYxcI1UVcBEl
ENkpmY9kuD50CEv6ORWfIkUdZ7It6BV6f4yXtgTxQtMOrqQhStqcu/AAqUZFwTEHYf478J7CNn1i
C1jUgQls/Hfi3bWriCJeOCpM8VoAVN7weeePYQUEAMle27XcTGYCi1YTEjT0y/kug1mKyH2ejqwY
N9mNz4g5nnoABj5da4kD5SvBm+eCk6A3SaRFgVMLNapKQr6p0ToWhdJPkkiTtH7jWTtFoLGCexdb
/Rwx0APFO5ascrEG0wef4FWiLIyiC5ZLaDlI+zpJKVwHbZSmqvdJ8skL6vJMmTsX8KeIM+jc8vQ1
A0VoT7UQ+75MupgS6rRf+sOG3pnSN3MvF2ufYl8jz5tFLvxpLjTPXCpfkZCwtIjSOpZi0+SZGFHe
QhUZGjMwtvK/DVYq8+uOv+xM0dNvi/Y7oxLHZIq/NpbICsTzNTZM1y+wy6DBLR3S7triuON+gzIv
IXqSm/3fb9WBgdG7ZNbeEg3yIuk9kkLLQ1KwbY6IijlJklncCwSpvIEf/H1p6NfxIVaInrOvT3+K
rSQ66XeRHQSaq5hZRVFfIg9qMIzCxQwip/oG8i0yQf1t0UPaazJW3KX8YMn5wZfrPLg9OV+ebiG9
PS5EA5Wm2xWD/+HfCI+ei6Mswb4Z0WMLEhZkfgpv5grAORtbh/kQjRpiLpBggpO+hLhmCeCr91Q4
D9t/y0vMo0xxpoii5ZJ15H5VcD/40EfNG66aARaclTzjC8imeL/rIQB6UMnBOwumor4cBi6SFeV2
zZlH5vbJzJccd0VYYbXIaiFET8dya4j+xyxVUGurkxjCjScIv53V5QZ6DDpBRC2FlOmC0ie6cP/d
SBFK0GP8xlC2lTEHlABMBS7QAxR4qIGgGXekGAOSnepG30jHSpIIchwZ8YpYTjD3HAJpa2AsuTRo
1er8E2pHIzKFCe9rRBYavo7ZpG4zf2tUH1ARqH+EMtmg2B/cBsprUKbZ95SQW8TJy9Vm4A89kUPn
vD626gS2GdUwcM7LTgXlDBB733o2R5iP+S/4qyqkVl5Di2Ahf833/WHlIa4wTD16MUqGf84z6let
8VBeetqjEC4hFwKM6aojtRlRx7BSI1zYULjrkobuBXfkDWjEBy2awBUp6ug5q4h85Z/PnzuOfqrp
sDcIf2wxHfYj3MEyD1oO8NWA0eo6zirlz71gpBw1odVVc6/quq+3TvTBc/KYz3VfazWx538CNCmJ
A+RJ9n6UoQPyY3sFmh1/XVwFaPoDIGu0ALKmTXJnXBs6n7qXIMO8jpy+Ow15mxxEgZsXMRGPogzq
KDbebp2vEbhraKSXAE/mI6h8h2zT7Z94RGweflL07UDMsAvnYpwmryb4Fjl0Hd9PfP2KKL0z23Du
SoFQz+XmHDRp8WWEtzEX8F8IP5eKglKk7nJqPbEFfsVdbKPjOEN0pXT/bWVLrGWlzV4Xi/EXLTcc
vEctQaL5CSAtt9qLhGWq9BjWMQ4Pil7cFvRN4u3F/gGiIJ/e6YD2wVPKqWgV2Lr0p4oUCrVLr/SB
S73AvH4lvfjtHCVpDUfnaQVNbRQPhhK/n2/3loSU4oANzkXcKcJuBT85Fq1NyLjBGgoU/uuPM2UX
MqLf5h0SJ3pSx+DLXcwl5wblJeKtTGq4P1Nq97fviBZVEW6ayHpbiAU6VE3z2q0fWenXnA60RiGA
YE5EaliU8Wo5oMus8gQ9yyQDBkDfAKUoP+YIYYGyRu6ZgpVM67ex9msyHYeEBtLcLK+FzT5DEJMT
UaWpwbahuoKc1N0kjKOm+jmRjNQ7Ns44sLHmQ946e6J5Cdk3Ikm1bQagewISGPdgHVb6s9sf1l/L
dNteDo45u/r/VyRs0IWrMIOr63SGS1Lwd1F+7wZess5LslIufZFQwa8OnMUBb+VIHcefHxt2OJHJ
YbX0ODXv2DNr+EkPPwYYTSTzrQc41iGUt4j0cK/sDiFqS8w5EEBqiasxzH2U3m3NEy6Shew9zNmW
DoC5Ea/tQ/jL57r1Eis+pEibmOx0KsUbI0k6CCybvJpgcGYGMLGVWBQJtJ0r7EgQTyRtZkE3Wagf
zjyEVKj5JQUJvmYy2tMBN49wfCK6ZcKNgIz7AwTo07RzHq0cEWQApWPOcbY0q8rPd9bHA+++Hbp/
0mCbcW4q4bLb0HXOVQKrOp/19R8aF92OI6hUdRYH23i3dLQcSzv6C4YxskwZtOqv/pu9lp7zHS2F
nwrNkT8F+MKbkJrDiZ2ehSFNrObPq9XPp//Z/MlYLN819qRMcXDWra/22eQfzV92GR0T3nsllK9+
QBdfKDIEuRs6IETeEyzEDlkP1JFrVjxKvM7cyIj8b9O3EKXZyYaspg7RQMHBz6DX9yryq2V32nTU
LMHx5Yt8Sm2HHy2rr9qLfLOUtZo4kULxWaMJnoXTUY5w2+/JIkpkAkHR5R6OFuiCXIOcA5Mm90XH
10VTfL0aEgUQBew6XuaWuEW22W22s8Tn1sTu+zJNXBoI1Kn3JJqXo5p1ObzjzmnSS2NCZK92goFy
JE0xkKd7FIq82CKpyhY/AvUulOi9xi11SmUft7W3G4YZxdWq600Kxv2rGqpiqILHhMQRzOLZpwEL
W2lSJrNMa2K+MkNCgTMOzDYwAXMKPlHWx0PgGNcQSfflExYl8SaCtHE5R+RfqwFzk6eJDIoZd+F9
cfUH5nXnSJ9yBWa1eqpQzM7CWaqloEQPGt9hXhOFJmGnZ1p7Oh3Yp4o8NGrcgRnnp4NMaWAtlGXv
BgE5co8mum2SlZ2jGoU94M7XlLUkWbaJSYXa0UssVpqFC+ssbGpkmel3Kz3797d872F+l3XZ3Zar
w6nUgOAW/T+F/I7qbQnvCOxhTiFQ3b5GmT4xv+GxBOE7mrmfqn0Ljh3oLzD4Md9XJ8OtCqlYxWJ9
1UEo1lrQRl1fzRFxHWIfxzQWsrQa8obncp2Qu8F3s6wOgj1F8vQaZjknSaiqiOJrKjdZtiIQ7iyN
awAs14C8Sk8Fj/lrOePpj/PPKB+/mTWBLr5wdzbFLZbH9WttTsM4uP3vsbRqGa3uVsBTgcwUVETl
Nt3DulS/o++hZGXLZyDhYPXDEQ/KcLrZQBftsGRqCrsyqhwnrwhZux9khLkub9rpJTWewSWkS0cH
pdp3iPwKKWby3dg8SS+f/lF7pfLs7g2mLKDnTJKJW4unTtmGpXWNYhSYoB8C5a44zTONLMr9sfC1
0TrkgAFsNwtttig6jiU9Xw1zxg+FwhjyX9Q3ZaeJoqLiOuCRwtFbkvBN0KcJ3oe2xgg9ZCo4vfLD
/iEGnRgTmk1wiX8ULhrADWG1cq0UkzCeXaZ4orwrhf4jVsHrWQrTwWN60ykhs8lJrOSykBuM0Oje
zOAe/WFhk6MzwbhR8pSVmzeS27qL2CPrWMBoHGpJq65PJFMCVoQZ0I8wYeJFxgC34eVdzcJFnQeq
zhOpusKi5PHVNPolT7JBkq6jncbA5DEJFU0W82e5QAKkd/wM7DQEsHVqjhqbExw7YibxBPf+hDLJ
kchsUQRZ9tAGkvZahWgTDKLz57pGUNYbiwEWIojIJyW2WpxGVUzyjyGbKqWomD64t1zh6hOjlZS5
12gHHAUMf9CMtMXhscQx8FmZRRFVeBrfLZ02lWP2TTJdqnfxUwfyPOMq097NXt3EHkJUPc4PIevf
URohp1KyhwQbDFooRGE/abi9wKC3qlyCq3M0qIEt9jpXbG4niUOpZYqJysKVezM26aOOkkQeFRE4
uZkRMJ6tPU3cdgx26qvrH+ITsdr2v9uUtqxDM4qJqy+qA857Z81jGilzhX6qiLewN4wfKw5XhbAt
pqF5ai4SB5V4FInlejBg1r05z9OpZ+8TLxvEtSUWZ9D6LyFhb8CDHLYkT5MAJ3Mw+fpTOSsHoVxy
7GxWGqhVLYXn0TlR6/9Pne1DUoG7S8UJnIsL2PXO3ON6he73F+ec3wVVSa5pmHE6vNZDNqMnZHBw
UXEj9/HZuXpzS+FNGVGtuxSTe64djdrMo2Ua4Fl7btKx8MoQLe3WqMIvOym5Kcs/fMPSQE3QGgDV
uu+ciNMeqNEq3giF5y3tVFaST3vkgC56HR5bNefKHjWT+Qf3d6Phd8Ae/45AhZtzbpE546YFU/8x
0/1mn6MccZes70TlFYDlou5eCGPW0jh01b3TQpkF/B3r4voYLVkMPkv2rCDXQHN9Oo7AFzCj9sOb
k04pG+rYdoKvm3FW9SklgJnP623iFXUZ7oY83SH5O1K6NHgVvD1crfaHmEE0RE4KO3JB/KA+YhVs
6jm6q+c/33XhEyCpvAYeKRQP7WpF5q6GIBLo0PjqPNCFlBYNfFzVlXAw/RUQR1E1zRMdNL+hna3V
2pPzAkH4g5nTBQOUTRjpmnzlenz2SHnpk8styScBgGDMZDVLIC+pikZwj9NiVe3e/KJqXZieP4E7
hTjEe5qhLSRGnzKyZ535mMb0bEc99B5CgdJt5dZCDro3KO0zkJodJPQDTg16/qO6VAg6j4+Wfqy1
ZGiqyfub0WgtoMmfzWZvTykMC0OhvMrVHQXvyYvvE9K0rY6Hmmobq0rZ6iNsggzpG9YXpWoyyqU3
DTILUKlIwn4Jspk1cSTOyPHr10noDAgj8eGDj/N5s9Wv65/plegvXEvZriz7Sk0zVYuElgrODHj5
RfKwV8XRQVlJcVexIzeKG1mHk4HKajOnq/2jgigNu1u7yN61IADKL9bJtHmiYLpZ9kGULiI1x9Al
LQvqNR7g/AFnrgCvYcPJWf51L/uwN8JiVlW4IzqWA4ooQnG4HEURi5l6tjI6AltHY7qgnKO/kmsh
gr5lr7L3FWVEMg646J/juD3Q3Urm+jxws6+4uIn69dqI+uAlYRn1/dOzICFMkQCQ07jxzLHu2ZOX
iAmdj9S/G+rJh5yeps4OWojMqT6TqX5k380N/25lWN5mFOJCSod9j2vjk7BtMDmqGSbbK2MNLQE8
Gkq8irnOw0rKnSxOzLSAOw8nX4ReDBHP4+WSuWis5fApqFlepJ7RT8Nf+bgCXupUhZuruBSWsEHY
VAKTWeyp1YTLC1sEU8exanVO8IgisDpiPFT7fsbf8E+ne5+JYN9qLUY3Yll3KXy8KG8cewyRFrCF
i3OZHx8IK1nt4D96d9wVAEY35UjltcOc1L+RR2tXqbUSc9okhivN5QcpUE0Qy0naWK6Xh8eMy0wQ
GzW75Pd0f9VMXDBp1/7hotdPIZ1WqUynX5qOUBNIwFfssm2NuSKJeaE45+Mje/8/W5R4Di8Xvy78
OyBV/joLzCv3NP4g5dH944sjOVL6UcSiFvfqKScF3BP6aOmbV+Rs/CM0QcqN9DkDxreJDEGSZhCU
86KmCJLC5TH57TkYAjitpKFLKaU0KzsNBRWiqisRwy2TPgzzpwGA5IlY2328kPtcq1YgJVtTVy72
fsJ2+8m3SI2T30GGdyQTkhGz9GcRbZdz85LJ/BrIXXAW/lR1qaFpmd4CaaHdOZcVp0X01cDEFzNt
CRbDHHJIA4DCCEhm+Oeow+ZEhz5KHUFO4Qbt4l2/Opb6Ukp+x3RUauR48PcfwzTwZ10jCVIIcYTP
DmR6aqHJFSVvHQDHnNdxViMcXkUMlbUjyXZOxaQGtMtMQ3pMnHmEZHFo9IDYV5fBvsBVE59RDoFq
Q3TcvTc44vVrJbCFCanAatwNS0XbnEAIsE96zr+BFKXW1tY+sOBgfjSGXHAmBBMTOf+FYNv3Vsd9
FBY1VVx1Fjroux1VlycSqSL4ksaWeGJpLyj93LrP71P0svzjgba6KyFck5YV3lMqw0LJAavNf/Ey
9xvoRVPCJ/WttwWRfRDc8RmBj6i18vx0b1maAj61di2ApqZ2HBSQycKS2IM96pq+wpU77E5AAgMv
OmHwDPwKzOWChbhsT6R/V46OLtiO6tw6xPfc97g+z0F958dJj4YFesogbDorcIJizu7XZbqCQ8kO
kvCp/5TyVxWVHuLS8RlKi6LAba7twYMCotsRETolIOJ/ZGy0qmGNmTxUcqc2XxGFJEAN5Y/b5e6e
hviau7G6uf4zCTEC75Sr/UbVSTKf1g7P7t7Gbdqm5MZg5XkU2smrcKl+2nlF1ScsCvoI2WWZ3JnK
+kjl/Y0nno3OB+N8onoiNsQ5wJWn/mAtSgZZpQ2XO/tbvdHYzhEEZCvw6Z/SnQEHrcENTYKb448h
98/BIk75f38jrdfnuQVLZzGgtolmYPZO153mWW6kRie/YhZiFYIcpMm/FQ9WQBimIfifjc/nVpdd
QiISgz+sjaMtlwDIzFkQ++r0I5SETSd4hLgwSZYg18+B3w2JMHCGBmZmQMC9Mx5DipkRcphNXE5R
8jbYlzhgzguAtGYrUXJzXhT+Bvtp2cZ6Pb8PTX0fcd7B9nQXPMS6koJ+SNUtT1eb2UiGoiLTNO8B
84LlkQfYmrOD1DDf3UzdHbp2vRb6XJTexsZiYJDjrMWt2PvMkE0OBuS8bI1RsvLUxDUrftgVevMf
4NJDSlRt0xBm2Ch8pHX2KqNvY4ATrIKNNxSxtoE5mMJkiLCEOotJh23qCj2qxQFhq6p5rVfwovAq
i3xLItocgBWQTOm/tMylchRjt6r09stvzn5sV4jQq6v7pY06nWLudj0eNvwW/MKtNV+qBzcAAiP3
V3DFKdvS5A7s0uxDSMcJByZYFC7GFw9ut7eokPw3Z0odZN86800c2j0qqNcDdOZ6mc3L7nw8muWa
K8MbIEOTCd502m/kuqBT+7OCBbsWDsIV1ogbiJI0v/tOp692HyNStpCFPhEwdPDbnqWScSpdrTt3
bavFmVBmq1HmYl1Vj6yO7JawDFb5H+djWHlGDGl0zimBd8QR5RYrOI9apK3XInQ+xwSuDjQmTfkk
6RuYJIqhf/Ihi1DQZ1/Dco+YuwJcY2ohFYEpatnCybQBe7ifmUxeYb12TONMB/cw5H4bkAjP4+Y/
grTMkKSJLN1PzOa29+9G/Osl481RMLv/hHzR5ezrhw8336cUm3SEJMThw6Njd9dzqw5tdESuf1lE
ohVxvai7qFwsXuLTpXo60Mml+YO06bopfFeeWbqwsliXmnKMlK3klnUjHKUnSB16TTEi0DyqSKWN
eIlfgeOmiPoLqhlqANWfnPOuWZFcqjj8vMwkfGmevwCiVPa86+DdsOGnNHpvGSS3iDP4ANcd30wd
5pOw8wFPCWan8rtWlI+w/d3dLWk3BVRDwhtWQ77rCIxJt5SsNSyuCDK06ItcAC5Sgy7Ivwt3GUyS
77NJ10G17icEBMr5JDk7TD/tCwqbxTZhWNsQaTiSlxZWeELvL4kmlHBLl1ltJtLGXyoAet/Ec0cQ
GQ1p5dDbK25FdTdfEV74zQ+MmmhMs7E3ti5XWBSrtRZZqrGs8uHWdZ5bdiExL9En55LlFOgd8rmR
3E75brrQi5Nx4a9So0wZqqQ+M01wI8nYj5SAAxbMmjPPwtpQcIntc4Tnj62Z1+PGwDeFRz47jLiV
L2+txouNIMGy0IliU38lp3PvzDb+G6FyCS28VMNyGqPXIffB7bLmw/IldSpKxC0uGv+SbG3j8mjU
Yk7bp1vnu9uLpqTnnas4QPfP+cHa3SZ9arQxvGjecGMrUBCXSDfFBEmO+NrS+QluxM5tNhmz2HPY
Ohn/JVyhfFgHpIMdkG61oFi1SsJzfcax9WA1eic8mbGx8IFEqJGBdSmBibFLIdy9r4iNIkrdnGph
FBLJT0bqOFxYexPLwlTHTBu6SPl1q6KfwbN9o6OYjU0GNm7aQsm6VBm9yz2V6swCZohItHPvfOSn
IjXTb+FK0P/vwASQFO2F4roIqkNzgwPDrj4yMB3owH2cttKPG+Es/zc0ny0C9W+vifcT6E4hLuVc
S8+rMjKI2fUrZLoQqU3uX/yvvnvLJIDKoqEBk2BWjPdSfgMf1Z0EoCybyazSd4a8ttXoSx3qJmnF
8SeM3V0/mCiqPJMpJMOWvYcWThqHE24nV121qve14bsFNCbMWQsWgZo4yqXfCL5BIuzrW7OxqipV
l3KaIC5+DdEucBuBRU6wCXmPnNSbg/mLTmj1OjVr+gDIcIQR69CoQ9q5Q7HD77gB792vA5TMISLh
93k0N7qqqzS6y5TMnLtUETIJIZ7FfMMCvwNEoU33hquryE8dhYer6e3c9i7/E107saQFrcz/h5Ae
nntSJfHl2JOEZ9ZLmTW3Epvli3uIV4kndVV9jNBRby9jSEhtk3qZeAb9IKPNVrNTTUlY/CQ7HeWM
sw2ON9Gi33sFii33KTZAn1Lv9zTe3f5uxk2WN0qPVX/qdtc3Xb5TWiTeRtxwCZ/dkd2kF4pG5pJS
66xWj6AUFip0F9yfbGNzdQrvKQ6G6uhvYULSDWh52zC/n5KokoAWBeF3BHF/+AtqB2mehOou9LD1
zRttnV7BCXYuEknncOLxeD4LrMfVE8RLH14lAMGbXUpfbQj9quK+tQ5wVUF86A87TNeueMCl5oPI
RE2UnFTpnUGbsgHUhDQDYMmRQ1w7kbymyK5hViDC9yli6hs8tOBQb5cWkHZ2xtBPpJRHeBnfhbBl
6DjWWbXEbgIJYeiwDDD570lqefxaCRrXRUiWDFvqz4gnSiC8kL8IPCklZEttYqEhSgYK9TiJmkxh
cX58YDyisBkUc9S3f5aj6Upshwk6fMVONIFstrN8taWIoMAP6OtcJou22WdAA86lffXPN9QjqYzn
p/ZQ7ye8f1i5Wf0H081ZiNYPmzLH6uLx6qmXQRszAmFjby6MJhqUORfl6D5lmgTzX6DH2uvcszY1
O/UUaexIwOtrlDI7qA/RZ314MtyW89taDKEE4kUuq7p/aIvw6mttjPBhos/2RlLie4JOx87TdUOS
NS/oWI8A1JYZcVOTpOoEGE5wxR3UJpMKzEmT4hwveCw07G/DnOZkQUa3rK2nPtnlyVhj+Hl4LPh3
WsSnr4c49/NyEbaqVgoQ+3sCz+SD6a1MTSK9cAkxHkMd0Y1HRQmlo7lBidcCGGkkEO1OX6HATNd1
f+80yGNNPU3/GkVnGvnkVhYzAARHNAb7t8zLYCf2wD6ypKYSNiJTypJ3vZOpArf3tIAsejeowNTH
hjzfDoUV598vDhWYSoTNLXA7SHSCg9iJr+cQfx0AvQahGS3w/66HkjYvMCNjDDMZm3XHir01qvra
YIU5GpFAMyVv2lhQ8j25D3P7wwI68LRZyNCdQ5+W5mbgq4Pm3SH2tWPrWyxePtmvy1WYKzRmhNgf
dCMrjZA1X9O/rT741aH27Vn4xDiG3pfpMjxelSO4hxCbJwqUPX6ix/DA3nmRPkEj2yCRPVULRw0i
dki7dUzqETv6sqZOb060m+NeYSxWn+8ZEfwt2HIHP+2SRBxWDobZ6E4q9CTj+kHD6K/VHKfTBpwx
auoTzFPQWca1lh6BeEBrxCDpXpRCR2LJ0Cy02QoO2EPOIKGUq0GiKxF5iqqc+TiYkqwu4zeYnRTG
xxovXQCZfcjfoqeLg45ep1J9pvFUG6GCDpHSuvdDqO68lfD3ASuWltqF7QqABPW66rNaU8f5Wlzr
e6F2Sm2am+gN6N98UbfqHQS9zs+UOsX3lWXE62qD4M8N9jaNuecphAZcxTSVp52UqxAVNa7PF2HJ
EZiyB4k9+7Q4dNzeBrMsHUWlQ32Z9Yerp1MQCudWXhQaHHMsca+2TiRstGWnhZHCRb9YK/5mMKs7
Rf91z5155Y1LM6RCxWUZM7c6hzyAIQE7XW7knPAUKO/Rix2sNzxU9hms2nZeXdlRyCQZO2FxtkdL
7XTNl+ixi753LG690sy4YcIYrXMTpFllosR+Fc84k5Nd3EMbmhch6IytBFao83VhT/ommtnk0/E8
+NHhy2ByHadkUkgZQNZ44xrcpT8lJLDjNewcw42a1n7yYhC+EAOqVcAdqdf7wrqKIMyQElJ0nmaM
OSNeQG0a8VePGWOy4XZtK/DMMURk1oiW5nfLGPgYurQLMW7jV98VQ6/v84ohyJyTwN3AWX+rYtDx
1P7TnsPqF4307Q5cLY9MhHdEUx/CTrg1LckFMYgg6ZRJnKUdCvePTjp3yhKuHPDKIkunsGrbVlkU
8rxjthE+1A50eu61CCOnZg6g8V+w7o3gvhMRAR581FUtWNerQ0qQteIuS6ttbl10msGYy+GwbKjx
KAdSRqmHS8Z+Pl5nB+yVSn12hlEBvbH20cRCdbcSMNB62/nDjeasSCNxA7NiQP/9Y2qr/iYMphv4
8aeLa+PGUoaQOSGLemt3HC+mhaLKBrqsysn2JMRU91I7uSUE2otNEPpIeoDgqycsONdoKpH+RIY+
pFWhbIURxTRvhhAo5fufSn7v2UBxUUqlwYXIvMn13n2Nuw1v14Jo+pwUDfSe3E7yIjjhOHw42/zm
cwBUqU1Rj9V4tiawZRPigDXyM0mba2PJ3oC0CEyTAsKpT7+d3Mk+tEgpRYpeL0g01XMgidFbIv1x
nL+n6E1Av9posz6chr7PKp5Y5l6mnw6zPZlCmQ4xfkYi8NSn81TG1Xc2Skq5EjWfF6LH6572cvP+
oHu/3I23FL8yn6KanZLcgz2pPETfs/V9E9iLyruiQ/LEnRy9iIkuO9oDKb8iDEu1PFF7fH/tE2OP
qB+GivnPfLOsConFo1hY2OrcpjxX0H8zUd/T54bNxmNHZWq2kd80B1Ze7aLzTVDqJE6N6KjEFu5G
HVF5XowkEGUpsCpFt+Dcd04CofeQZipdQYUMf/U9eHjZse/mv7jYp7fELsl8U0p94ZI4NjTVjaTD
qAjXAgSG0rj4fz8IfYNZ83AH2f/D8d+mu5NfnicvfpypvyijI0tAIDmkUKrTgW9gwmsm9VyVao8F
8+ymIcTAYm6TFow35uvhy3EDXZ7KFdEUt/0nHok7H6LZwvbdvWTaDDg088icJYIhP6KwPKKAfGBN
ULoie0ZC745nnoSoA7oP8D850jv0w+8hk/L4SWp5di5GaQrpoo/Yvae+cKvh8ZX4MNGVu0S2Y0pG
4EGVEpn/BLp0NuySpUS+Yi7m/KaGAEY0TLkyFm8NnHBV7t6lMKX4Hoz1khZauM8CA3oftWcxPDZ9
jyN0eMICM0B3xnlQSmMSDpEPzW/WYKh7wWNG7zGoce0dyiJvhAfQoU3OBXj+yvkBOkoKaCRTjYVe
NAxYiNUHkzfF6o8b/cXO4IM/7l+sDgUvaKGgdQvvRCdyML0/I7D7aVSIAphynmNNxiosv696ZIum
PvfVI16l+PmAa7UlEfIINSK9y99lPbAKr/ogtWEb+7Rk66bqRUBi3nKzNGB8zHLmyNKDPjO9mdQC
Z/hqWkbdd4mXlZw3fuwmT++f2IU9u9VsvPU1xCfve/LX/UcPi2DAl/F5Q7BlDntV/buZ1t+5uuwE
3VdWDOLmB2AON3+FG/haIKBSpCu5gwbgiJtNqGTznwBHvxue6epRdjS6CpmEKi1CeQAV6eUajli8
E0DSTbQMw95icQt1VpyGU2Ae3iPocDETipJafGL3cj+D+EH+qr2YBBaLwSXnGqzI14bbuDRdC+8K
zu2J5YGKYbkNmBFDkxyXWiBswik5uvhrEEnnaImbzt3g6gKgjjxRJzZnbv1JbIG3puz9Sl1Vc4Hc
jW+1PGcD4rAvAS61PhrIrS2ErkHbVRLdtxY2DIP7TfHu/kTwGmTKG2EqwDtim7Vf2ImkBsvaIKL2
iV7D0efWk1sHRjlR5Uel7x/hhP5OYYrkNz2tbRh8hKQxOD+7A9Zyc6hLb01qXDuO7JpoH5whXJBV
EtIZmyvzxGWK3x3Hj0m1rlL7hVFO/lp4C68G1Jpy6jcjV9ZUJ7c30pFXO32W+fdBxeQT81VN8q22
9p2l5hIzr3fGp8doqwNRhCdDA86B2HIQceDVFGn+2SCRIqqcM9nPJJ7ttaKg1e670Xb71dXb3AjS
cd8eiIXxb7R/vAR37uxuSmoHBZScBIRf4Pxta1qgBSqGseQTnq+2Jqx09ZUFq4ZDSyhCttTn+PLV
mARUTP7MoDXoh7vBAwhsSuNstjYhTW6pUTRs21IdjWgoS2OLLvlCFSQefeyi6g2Qa2Ii2L5LFDzp
aMFfoOMjqRhJNUfDpO2gC+rgmP0hh9tTJy8RsZu2WD7KnXg5ONW6+6ASVRghhTnS0HgYvaQSvM9a
vgMW71bJ5UAUCnJviPQQo96liR8AaiECaum5abkLRRYtgGmKKT5gAJwnqAHjjNe7J1zZWZqAkS7K
gz+wqBpiq3kNjRr9V3XZjk3A4oeEn+kbqE1xxYLagqChbHkRcdLtJRgcP7gdi57E4UI40qiEppE/
nBRGfutbCEBVelWtUMacltsOTnjsMhbt1btUjR+fabwxphb2sIGIWXAC4N1NsyiTRjBlQLT+RoZB
ruci7nWRL/zeaXcaxWvHkp28ONHk81L/3vIAuia4DF893xeayzy9HfyJW3PXRAR+F7ZMIheXKq21
TUXrOwDQejEyaNMa9aABDgEU1Hn3kzEZ340WZtNOvXScKc34qLQQz9FXCcXZ2qznXXq8DsuuRrL6
Ynfki1xfwu8OfCFORl4xWPE/ChG5jiFwezPAuq0QWeKRZTMWgPG7GGSiOiyGRzQXwyznc1o3h/Eb
5/KW/nDYwYp8BKiX9+Xk+EMuwz8bZr3WjmESumtk17qr/E5jpeH6qX+9SBOTHjsJanu1tuX5Ahuq
S6IaUhMllaUI0zdfRPvkcx/YCUK5Q+g5cjL/9ikmFdF71MsF3A1SG7aNWJIAsgqGCnVhkzNQoTBN
Ephkjqb6jjSV5Dk2be7xUh/9umZdUynlB0mlyOh/XcvCsGfTLundBbJ6zBe29M4lAO4we8/68vOi
GJScP2u2cRqKMWuXVbBk6r+3X63oXE1mI6J2G01KAJhUAX1QKfYkmxbRbxqwXkJ5wuzy4dwuZZmc
GpBNioZg9IvdzP+lLoJ1LUmouaW9HA9DmrRrIxryoJCZjVUn06NlDZUcX0N/gGSdyHgIt59j73Ft
8lqAlHa94+HPzaDKeomeikxxRC7IwXdYq8mHZ7ODxubTFYZ1qR5Egm61L8lDRMJSzoyHwc+7R21u
7gvjJflWN9p3fMsLmfYAxdjFn8i1Qg+pcfy25K4HWvAkqPuJAG9gMn+Jeh2baAGHCfQagYz+UCwl
cN4CBpuYIKubvmscpJMn86LLgdt3NuAYuMcEqZEEZxmhLCGP38J+L8iX7IqJX3QB+OpfuwyFET74
WKhXpNdADCIeczx48ILUclhHzE4O/zkIB9I7HyqqRxn3KiXJyblGojzLI31TBjVH1rWbfMzRGC7E
gvSYNhKaKGvBXD6KndfIccUKVMvN9LewaOqJSSLNgBY9ppbDt9ndhyRpTfSRdJ8DanPiO3TrBfhK
FiupJEyEMhN117XRyiGV03mCCZv8A7Xhd1uabVv3xotPi8xkYSsQVXMRQBUjaAZuuxEMNmxNVTly
8g3auLC8pp5B/5b6XRqwcpZaQRZn4TzYc1meNluzgOQeB2nAQr7Pmp6Apy0jz1+YfB9KkwoWqDHR
ioPCxJXGbgCJuio+rMeN9/dm0SmBcJy6sZXKibgOhQAgBa8pQPNSWjw2jQYnnl2lFdxjv37DY6TK
a63aa9ZseI8Tp0VgUi46eYQ761E76+RvhrHC5pLdSRrtvG29zccQCls27vcvejKw5bHjn4GkbL6s
VQ9AWIcLOFhI4FQI8kT/3naS7QExA561fdbMiZQLEk231dObIrJe36H2vCYXYkmqr6uPOfqgs2gd
SxG8qIUFw86d2EHiaGFE7u0XshNhh4l88QnSa7z1mA1/kITR4XL1HM/u4MifCrwgxIgGWRhw+SVn
mGcoZZPB7aQqsCLTGzVzaqNSlG3eBY0Jzs4uLq2MLTm1XyDXb2fNqSlFlGa5uwTRoEvYf6d0RZwC
HGenobb2d+9hdQEyrpTltnvOi8LI0rjO578G3jzX0KybkPRmezYdc9ZqTA1ggX3InZLKnItxMSk7
KVqRd2SU5rQ5jAlt3dMMYPw7jNmlU964UUV2CAKa7+9/Df0mh0VLPTNJd2rCJN8a7L/albnR1Z0J
rwRZJ8fTAod/7pM6pEhJOV/CCQ7E9S+T2h/2opazuRRrXXf4cTn6WIMyubztJ+84vYk7tpNi/Z5S
Os9F4WBGmwokWqVBKt7ABir1+W0DIxxWXzyexq4T2LJuEsTaAz3mDsCsg74asmgORDR2U+JwAkoM
nlorp0N64jeMuvdfcLSV77uzouirTHX5U7F4xXXINE/6oCKu9u9+e1i0SqeitZRzCu9xf+LrOzVX
EgHGx/GseguB12S6KoLfUwvs8SncNUlrl7gsQJVfM0K4jm5liXFAOEpWuuzYGOcxk6nUqepuew/H
TAcndU2V9MiXRRGs/2aCtSMEWsg0/Xdend0pNZcn2TQq8xjYci5zvJ64UY5/k8aBvLne46JLIq3z
Rj2o2JuHjuYn8dsdjZoel32LEH/rEd8LuXtmjLcpeote2MlJxxUGJlDQleS81uZyPwBFdlWgD3NS
j6va+AI9Kj4IKjvbOKOKbqdghdtO8GdL4E4+NG87Z+3w4pOn207h/1VmMkpUzmiwLD7ON7srWdnh
Mu/ar39TvkBXjxsBRmMFCkxMyNTCyhJwHkSaXgwevxPqp+qZ74tPZPxBSCkePuoeQYPzfZ3hKlGD
Tmw7fgfMoE0LZlL7euColzk54Rm57Lkdd9txdOACy0kinp5nwrqdN9x3z+FnHsmEge2796OcVCF7
+MpP+DJE0YbsCH1pF0Uu6jCN9JhEQa0H+POYXDK18nxsXt/vLLARCro6apv6njCxb4qW1ROpzvcD
cFDZW28/uEHoR6vIEOa9z7vllV3DggkfvsTJ/5FJ0PsOX9aoY6iLSqBCzS143/XzmtTFci57GXIi
efHeS2ptXkg+mtNot4vAK7Bw/EkKhiN+OUNggaT3iNRIHHSRS/9mxJ3l824oZtApXUiUHCMO0G1V
YeD9iDlWMDUiJirbYNBIplQKA7lZwGB0jacPwNS4eDucaeZhq1tjmJ1nKaHV880FF/FeRmJ1hrWy
wsHb7JLEICFa+iLIa1PWT3o9JjCqcC+Arux789CIFtzsH2ukDI3HXtTfg1Vh3ITsCleeUy5iPZlQ
+iEt482t+7E7mAle3vD2Y0e+dKvWqhVjnEbZG+r8YbqsBspC/CwWnJLL6jCRZLMULeSUVsNTscuS
/Ml+jmBh0pmuwG86OlIJT+2y65A4RuLwhwdRORjtChiyuJsW7SiZ0TALZeReoeqUsRnanpdyNp2k
perJk1rrR57J8KosCeytlMvG4QpNnlfcxALQyZ4fdB17ZoftnKJqSMQgTr29mRtSQsuVNGU/DOVE
/rMYfVRWKNX1qERoxaWQEw4+Ra6SNVm+IuisfXYpMuQssQb4dOaWo+/zLg3Z/x7SgpQ8aY3A49YZ
MWOL+Q4hdeGT/GCAM7NPOWXvKr9HR84bZwz8lyYafpBttfjlUKMXH5RTcnzWDYnHyBgY2TXXt+pD
d5pX5pTIBQdsPAvViOHd/Fjdl4Xi21ri6dhFOOONyY/oMQ0F7MCgsCw7E85WYCVduh6mDHCvye51
eQDnzeqt54fdQJRyBkqbSfBJTNZDBMY3SVzkx8x2xN2AjaEcBtReGRnpEkBLDOaFvIv+rxuziTXw
6g/fyHp4zpD3BM4AjoFUdHQP4Z2pg2ML1LiuOZlEgbkeHmslgXSwfqaLCFIpzza/CFfwUporDNxG
QBIPGFm1IXmUQT5mcJdRaN6vWPwxlcnSl43lS8nLvPrHYtsZngyXImsBwl9RtKmyhwyo2OezJWNF
KRyqjZHJs3tjuwOmBYCnqvfy0aj9U+342QpbGniLqFz60zXkWs8AjJEDbrwbIh+mBTCYdIR4ftrX
hL1YdjsBYhoXjHcSvHMSlsPaLCClBVU76yYI+4pQ7SN3QNbP9mikDrifGclqebKSypaeyHPpkRRK
T/wNN4t2KQ6AgmitFwdNAod7kfHIzKpl2WiwURtH47XUwatF9qEYbH1DLruVFBRiet1S1RjnXFzZ
GKWpwAAQvpR39XE4WCod2pgUewn3AK8LTBTqFTMASzKx5frojExGb8pcnPXVTleOcVnMqQpS8Hba
FU3CIHea8sFjMPb/cH0S3YT5xqlJX4o4YsTOE7II47zrkXsnr9ckZzRjVRCboxM+ZayGsQMxac09
p8pTQa3O1phDjDUnc6X1CcmTruM7DvxJqwJpVMZt3PASOgp57zh5R/JqCq4Ru3f9xzDbQ47oIONu
zQW6tBDpolT+s/DnqiVtNYXtxUzm7bzqsETIFvDCXU8iEXju2nBTJXE+SnF2uk8CtxIsAoiU2HLv
zFkb0Od8OAZPqIqH2hreEBumQdnToRuq3p72WsWGOIb2qZplFTVEvG9bmPElA9hXzvm0BHE4KCOx
Avw8CqktZJnPUtST/Zjwe8fvXLAi7ic2jZXIF5qbOpVBbX4AmecQkmeYF5dLgbqte0UqY41aDmJ4
lltQa5EStOAPHlnOsF1mJKJ3/cFXOdgMR0OiLhQPZHRU6YaQUEEHU+gJNbzP4k4HKUL5HR3OeWVJ
dyH+tBKPZDtvhNlf8mcbLVpBnLUkPsyaD1KMZRQJJIq6i55+XYrLlfA8EUbYB+SQWd+/DjdWhuUU
MkwRgfEqK7Z4Zmq6eiCQUccFXfvuK39yjooDyblym2dgsyaJrFCk6wT6WVJnqUjxMvm9/h/SY47i
CBStzi5SBR844RL0oCzzl+9sKshAYF/gE2AAt04RtAarcpvIVwQFB7ygFxaqnMAqc6eBnFZ1Yi0K
x07/lvVz9igMOpOcU9PZZUd6aqVvg+NfMy0NF6seLD7kB72Pd+0bMqRCSVt7kGdSzhmnLvarvz/8
Wh6yylcFHypbPbfAn52bXwZzji5TGIrjsTrSgY9iz7rUjo9F0dGq4ci9JfJWaReLQf2tIUNEt1bw
9cK6X4s8RdT9m5at920nDRndx4jyN2I0R87/zYrdSIBBPl0cZ+WHv5Pu7btmDcGnwU4eSKgd9rBu
CiZvoMw6rGXJamMvi7ZC9DE2U6sz0O4VdBYgO/Jmopc99TYxE1aR4lH0PSAKqKQf5wCrb+y9rUH4
Fa7GwC4raz+ZPcl1lDp1MmZP2c18HWZcNGW/nkMdeCR4G1jUw1wyxnaAPmQ/dEMSQ8EXq3SJPcyD
n55uqHy09q9gAeXrKIyOzJbhD96IoGeQbL8DtGl9/XANXw78qNq6kFQ6iQ90WRX1oPSnAgpOUhTr
S5i7f1fQm61NaUvexA21ZJhgIxKyDqqXisAlQoyp30rB0I//FwcnJvVvw9XdxhWX42seaRwWKDKZ
46oQm1dUdJUyry7sOqMo4fY6v8cL72++dsYp1Yan7JHvX2rzltjie1RiF/wWGHpKpJmkf2Jc82DR
vG3RMHNzzJ7TZkzG/fSdP7m8JhO7AGx4ZuRHiKPy6KZKES26KTfMp9hxfdShJNeTmE6m7Iuh/Az2
V8wuc6HuByIVGwNIQX7vupoHOhbMT1qkYtSXgymmIl9AjgSanhwgAvbJ50LK5VcncrHhmMbh/ds5
i7fLNAGprausc57EVMtckMvneopH/05gMgwYRISyqEeD+oK62xfg8D6VedwGyEBsOq25QbAAzR5J
ndHQo9Fchcj04qWKqh+o5dqWKUCw2INrwqkgT3XIgTa2tBMHa7jRIOn6LvApyrazkdMyvmABo3RB
lptCBKnpsg3SKVZ62v7Wy7PbNusXSd5VGKheF/iIHkkp21a/UBxWTmi5pGsOyzuMDECcj7Ed/ShQ
/PIsYit+fcYA2Dye7M+rKC6QmJh4iB5LZnKoq9hH4WQtQN5sVPuOzD1dQg57XJQ9Wfr72LatW+G/
LlgtFXYEPmCvHLmCxh8JdWu7CgcTFbijoQEtiH2zsSUOaelnB2py5AaTm1Jz3DRQqRke7I/0O7gt
7yoMVHp7xK/4tjaCcV52OAaGCJwNHJNqIBZ82am/U7FExJ3nHb23qziHUJCFZ4iss3SoQbbwmv1A
uPG8mt+dI/OG5o++J7Xt10uQi2B6pi/XjMVv6Lxx/choND9VJOGBrzZUJBJhNhqRbF5dYHLPF2zJ
1AV+lWwfMofn3wcoDZBuYrJyVC/XeP5h78yBJjHqy6cv94DSUIr3l7KvVmHeZ/EE3VzAYCwlp3mq
pn9Y4Y8X07TCSS0cinJFjYeLiuVf2F31NUfKdZtgiZZTwH7VKGferOAcG3DAHIkSdT5Iv1op/Jdu
Y8awIrt78r3U/TiSRcSTLRImMU6O4JrOZXCEqf+qREJvgBhajHhtymT1UdeDNyBKjhmnh+LrnemB
OT9Agr4zWe+oJPg6JWOVXXp96YRaLFGdSYJ9JBLMJpauvmvJb55bMtBNrKGFTPA4P48lUCNW9k0e
nPLXddoK+nPmG3zmrStYpnQKrXQw1TzGNKPFG3trvUZLlMxEXyjol76hObWvGYI1PXr/9/EV789p
BU6V0ZnZ9nzMuTiWMBbgD29YUnVtkUU0GLcoqiyliPPKN2CouzCRr6SKGPnpkQ4Q819TmuBC+Scq
zCoD+V+tKWqjNvEmhe45m6975HAxZnOoi9coS9375u8/5Tr9iB3EW03/tHc1uWcJmjIy4TQqpv4U
XqMgz70ooHXVoC5eHTatSVp3C6f3PReFQic4eNvZmPpqbPUeVObwcYz3TqONMAMlPpi8v4NVg0Bj
gdkLgLBiGHGWVYS7J4N0nvPiywoFGJ5xGnRhH6dwek0fy9odwO6iW3uH50mUAMNU/sBBaAQr7zFg
DzzL2WaNSmwPhEXI92k8iZL7J9JC6+KseGqxM0eZr9HBeo8carJv3bKJQHRnzZjN5tMAGqEqPBQh
ZV9eyaQfGDKy5haEqDjpmqxc9t3BwGIMHGx4xoKjBde45WAF6hxjyipPsJk1+K481K00jc0pzLhI
bnWS1mVrK1ezFiT76wzDootD47HI7+BFwMRgk/0vx5MSZcj6Kl4WgDV6fAdj7rF0dfeek7v3ORXh
lcMoy3656eFnr9YTXkJ8hbN03DG59QL5xdQGEKtRK/4iUKsTzJme6jdnNDJbKweYXReNnujt5JNu
ax7n9kKTQuhLQSxtddRrg6wL1VBgUs3Kr3FXcToCTRHCeyeO8K967JGwwBjEi2QK9PikqAmnAOMf
rPl2lJ6XJy3FPVzkq/+uqVELe8vBh9NUNm4YgF7DJYADe5b/e40TFCkjEsk3O/GaLxuhXoLtHjbK
CKiP7GZVTSdZ58LMcnXH7kiNZHgSxPudy2rZGQhCfBPsgCkwjPugtQ7DWYBo6ovC38o1kpdT1Nnf
aFGDHGU9uMcrsWvUJFahjAkOxOG5LE5nQxOb06VrOvSzUuPS1yAkoxHUES1tmKZbtXBUwYsbdmEk
9itPmUCrFbmRUcJz0oD5jSr6G39C2p6izfpw0sh+StlhJE1JRmkynkwHL6v5NIti6Y03tIYyaBko
xPn9N540K71cwY9vj9p6xpbLBTnFqQhC9HpTK8SqHXcpWvBr29vQ/bJaociKZ/iSnl1KQX4c0qQV
8c4YfYIUJu5YITsdFsuuLO4bjH97Tp77TNdaSioPhb/EZ2ynnyv21U0/wpVD3meuStkTa048w7n1
ouhqoHe0mYx/n3I1cIcGUtmxHFM/Btj2eElHimuXEZ2WeP9pY2OJFUcHbsx72z2uX6U+utfYRduh
Fh0sDZSAfCljoZW2RgEw1uPIl1gLu/Wj+/ZV7b/MRxj3fpPgTCCaOHyPBrbmzqLsHD0yesdjxl5e
SfLUN49neWzSwr8LI5yjhY3jK6gGXQP2sNsdF8IlcMrsd2t1Q7CXT2nMLlag1yYzPLEc3sylmF5i
32lZ8cwPjPtc4yLHKg9CgJaphCP/02QbOyV3EX8s9AXLEHJ/QAY88PCMFDE34kRVV8owtcCgF222
hKgiNhW0wk6jvIuPWRW0d3ayCM/RkXScHX95N8CKXj00+Np7fK8EKaVNUgtH3m2jIF6ANVkI5Fo4
NGCFQLB88JnAAnwC8n+SPGNFlWS9kfx6HC77VMzrhUWNdPnV0y/SOM0WnKFHhIWNpORWGCwiKGv2
GHyD4HGvSKWW87GVQ8mjUQazCx31cZB/PafMxYzJTrOHia1MrU9NC4WolJ6sSLT9YG4cUuN/dvZN
6Doqs4eRGXgggB1PzQ7lOrZUigDtUIygLfonm0tXOwKNP4IKB+kqsQ5B0r+ww1sRyRPGFb2zc91i
xRuPOXLKU+HEegznRPWrKyXnmCmhlHaTS4W3kM+aQGJDXAdeoFPQzt6zTSYqYYam6douanyaFonv
ljunqO4G6qTala5+dDbFxOEJhVpGCwYPLPnJfUJD9UJmSfJ2qRrHitYVldEWZ+XAjFXG/DY+uhl5
3ldZ2FptFSC/2KyfA2DtAmkp6SWLLBDbo+Oh7wFscn0noV/4lCqtR5OgwCTIC4QiWEy0/TvSST4b
2KBP8Wu+vwX9mrppslp29wBTtF6dJYGf0m/0Om4wXYnacFUawvYFrXwWwq/muWPRuj5smxCRo+dm
niMQBgt+FX5N9WvzzO2PzmcHV2wSLlpBPMpa5zV2xt7+w3kWxYxg6kNGcq6k8fvm1xem5cys01/l
1FRdq8XXQzd8+OTAVaxSS314DpJJPTGn/Q7VVdiPZcv8cDqcGZGsCy+XoG08jekuHKfIWHwuHY7d
hif0fq0RSG+eIO0RFCrctNqLHnv4Bg9Kp+ELejddjXw9VXIYb6O1jHbtkdxUrVdXbFqVffHgOccG
B8gN22Md9i9ZILtW4ns7c3d+bIWjPj9Cyk0E9Fjt0aoXYd3SaDX0a5g3xvd1B0IZd3/19ClaJ7rO
5odmgv7UInm7+reTaajOJAOPuZTQvqqFtcFEIWENCQvcjgJ7TMiEZFPDI7gS9V4DoiW8pXmGGu73
MkmQi19OQfMSk8TL8z2zNdrs/qJP+mOfTQmbB0trcXU8KDw/bfzIh+Jo5qaVJzWLX20TP1s9o12o
gco0U+Ha+MZTwifQ0KAJAo/mO9kUYjR0a4jxd/tEukx9c3VGdkLbO5XN3jN49AcngLgb7vJ2Vd8l
1mAyvm6cA81xMsgOT69x3QiW6Tp2Hu/hWJO8GuwHU6pZisGx2FW+LCx5Id6FHmHJC4t3MkC1ALLH
u6g98dYNWVMmUiWK0y9QiYoBXFiSl0fGdyB84RjnnB1mJKXJTHQTmhszI3IJhfh5g7Z8k+9s5dk7
lJ/Ph89kdHGVguj89S8UHKs+aJKE/bScun+Fh2L44fO3g9hl+6izgE454bcY0GIJ2occdg2ofsNp
Epg1VxPBPvPXcwt7stSv8QBR2z1v46yJptsXP2KaGp4foI4wY7wSCa8Cfq6zEH8Pb1wHWNFgwFH7
7dw0103seH+KR5lR1X71Rn+O85c885MT9nuj4zWNkVZy4GRz0QwnLakvCZZk0NjVScHy1GG5sKHk
vjX9Eqe/1Mlz1VC1oh02TtPjy+7t93VtFYIiXwOlGaWFAIy0UVIwlAdy4KbeWyXMXFWNDz14wHHy
uGOR3RRkxIMBETWnZwdHquSAAhFg1YRMS05l8fU+wZUHPa9IsY15/TKQT5SunQoUaKt8WH9aacyh
Dbsb8YFshYZhJE71ngEU6k3B+tWBf5ZrbmGDf08vl0qmy0ShkahU8lQKBUA/yHf2QtJp9b9YoT0H
ZIcQgCBcd/3Zdxcu/nIIfB425aT3DZdA9jLg09l7nb2RwqOcO9+BGBDok+LPgfa2aagUAFPikYUY
YXwuOHgF0I06svsQEWvuczRELK1xO4ngPtP8zAzLh/n2F2sSrHvTnTJjXNyIHzapmV0svuRNNFk6
yHODdz7AASOoUXywojZ2I3LOraQWIp7UJV23VazPvdwLyZfMSGkeJ619JMDHa0SJPua3uzHF7MXf
bGsgYXrBsEx5n5Q9HuOuvE66eQZr1gF/3xbDqhy5FHGmBNJXGJWmQt5OwbD/ZfmeqTEYVwIRvJTl
JGsvLosx7cwb/lCdnXnR8xDuHfhbdj69pW0RhplKaneGiHmSgJSaDvJciq4mp5uT/mKRCsHTAZUZ
J83MDcgnxaej/DJHLrhcfUGGID+Rc0/D3SFC7pSkd36lt7kmO+Hhvko4tN7pE/6OgyOYwsk8hiru
YvLC2fHqfwnEL2XGFlEtYIolNp5pnPCEHjXMBv4oL5uEhUBWOakMrzTpfz2itBtO9kkdvRb/cuXa
e55X6XUM4yzvHUPvK9gnYCaGpX7sGkJ0/xOAizjsR3gOQ8B4Rgm0NKDJnCv7bWc/a2lp7MJ9Um6I
+FoRbNKT9raipEfIaVqmT6IWsBZtz4EVTwkVb1hpVsW8NL01+QjIVG9vIU5CXTfJ5G037IiLcUuW
bSStVAxQDTu+ANuJLls0+6AGT9++yLg8s4sBu8p08xJ0SsbdjlrQCgUaeFemGjtyURjyQ3HPFIY2
SIkd1D2IlgGTgebSoxnCRwDG3045vlLEl4rp280oYBYKiLUnGppBGKKiulBi2+xfPhzqvIWi0X/R
1HOakMl6PdNpibaUAbDMwqXntl+UXJVV+HyljOeRU9mf2os90WdHHYtbWmRviX0002qMtHJ9be4m
G5b25BL2MOOGQL5R3UGQzOre2/CvU0GdBtM2OCxckF5i0xwLyKktJ1PFo0TkLHb9Xt6oStpa+7Q4
Uh4NXUqHbXtu4715bnF3oLvC01QeRntN1gBbe7aGKMPZ6dzo0efZ7cLJT0owmNbvZko/OpAu26hG
Fl6ciSWEyQk7t4j+RELGs49K5RJCxGBp5dFVICAu1cNsNp03zrfQjsW82YkRhppVkbpTf8Luujja
0thtKaBvsYoCzKhm5D/4EED1/fFs4Uu2LFV7r5Yvpd5c3H3T8yCFt43sFDGuTcYE5OcXKS8xTWLk
4ok0Sd7cjhILbPyTWOLvgd9Iu18PQkKw1bh6xV9X8VzWz/WDdWArVmVvSPwgNyuPV6FU8mnVGUkJ
0n/REh0lFyL/zVtFVBwu/ap5KYF3OHxhFLr3BRmv/thb+rgSp8OKTLv1H+wD52BjRP/oB7u5Kqgs
Bgz0XmnpV9iZYqYfK/ysbpLbC/ymHBs3nBVlaY4uDAnHaxqftSX8znlY6a094HrhUh9ijX6EUhlE
27g21WnEoCo+b8/sv7nDpzOoIRiTRKKAyTu5oh01aVRdeDah0evyF/1arI0lnbb0W0hYvaPAdQk6
FXa+2dn2StLy32v4efJRspbd1d/RCOBL1ghhWG7ZrIJ3ameRAHUpoD+Tw5rgqUWub35cj1CuDrgs
34PJQMv5ciFCQuPL/kqtD2JCh6EXYJolrXvsTxU3ASjDYK1tdWi6yUATaRZK3fPVNtGH23yX/R7m
LZM6uHnzm/EDZHY3vwKpqwKocsshBARMF7VMEckPg/ynOd4ks2xQ0Fe+miGQEKKRmRsRAR9bYe50
4G637jt/y6/D0ZJvbIqpbF7psZiV6nEvwAJ3JG6vmtG5HBWQ+oAjmlECbyM2mny94jUuU+npzT4Z
U08aPaurGDOJ650wAPWeLzGq/luoV1Qe3FmtGTxTQc1S4kfmMO+diu58R7VrlrzI0Ur08BjkK3ZA
FOXSDczHayPK5ARUVbFRQ8JiAEgbBAatsdDLMv7agTfnc0nvi2vyr/zK4ozxxWEJ2b3DDn3IV6IF
3155vVPJ72fIFLe9z9y4pYsGM9TmMPV/cudx3FTXjjUjWqaBIOmj7Usb7SGaAGi94ImlBwX+A2se
pd7YQwQYBqfNKJHTaTSuCybAp1UZWIdUdjS44jTe3vNjTLkUW2gbznUF5/0v2Zhj1ydZsYrFhocQ
NYnxGFa+4rc/Ppcs6717lgmowirChxZj/Z30M4A70Wl6+jm5Y6gVzHBoCSf/VYccEMJYLR2eNwpt
lr7a5EVW9HNcF5Scg07VewxmlKevGVggiDOWRItzciiLFAT1B24XqPE9sD9LOYN/A9yww/wfVoDn
nu7RgOUnAXtcVT6Qu2mnaEhIFMHemxSN8y7v1A49Tk3zGPOZpBCZZUrpOjGGELQdHr0yh2s/oq/s
yeIsRqvAau9IIBZnh23kzFHEKsNrV7g6dGQ0CZLobfRS4xoVZDVUjRXQmfY4hj23AFS3hVliVCQv
6GEtuTYlbBnWY1E7rrzsW4gjiXrzTlBM+FXPxWyaBLPct9w3sUxPHFSSPjdtsmMqXUuehjwBNXHG
I39mmpdwL4Y/FODXTpMnOXjzeVur3QhCj8/twf7mM/rWmEhPYYks7deDhiWYKvGoenhykSUZHruy
TxYqvqJuUovRuISoWlv028VhMcSOaiYdpi1Z7bP+Y9pojRWPOxz8rh76XS3MHjQ6zAEFg86bfWZy
LwjTI8bMhJf07OuTiRF+07qm1U1KZo9GEYx/s+mYacozExuwO+hVY+6m1RzZtrAsjwPGg9JntBmW
onzfH3KWU42uV3uX9TAXbql4iAvyebptM6t08ldYoyQssgvHtE4Z2gn+HoVDlvvnleMsNu1Cj16B
7UP0lDzzSfP/RpRcEAdtGXAn48VccndzoQ+VRzuVFYO6c2j6gxoqhRjbX8zCDWPGSoD5I3Xr6Y/G
3rUbE9kXBr9cI6ibF+uTe1TtJEesetjwL7FaHfx2HIs56XILZZuqoJOLUUSN6OJZri/dvE6l7DDX
gEV3E/g38rlYlHnugGziDm+jOhQN22bd8RQdBymySV7nuioanokarY51iuh9vxIMWVWggZ9hqOE8
7sWz0CrmBY34QcXuQC77CPaGF+xe5Gu2uYuk4gd4L40T0oX1nobnjyMQR3uo79O2yftJRMs2HARt
dW6AQjHURT6vQniRDo3ykxgDUp3agOv55h60goxDLXcET6tgxttTL5MJBZQhKUHCehkCElQbfmQw
gl/RpS2LEVQByc/sj0z03M/t0bdR0Xx5OHDmalDohLrtpWGzQ6MYhrPT/qXjvhvrEN6oJrBJCL2t
W8FcQxoZ+gmcbI8nOtESoaKcYyAE8O0+l2xazvgftHl7Z9NnVkPw0cv9cmd7XSrDRjPhRPHxfCd1
v8RIf+VVDd6YTGQYd+ND/oh3kJf2EvtTuh5IoKOd0+rNOjbUo54AUsU3UvzQuEA461cVQEX0hNG3
Pwi/V6D6bK4/FGeDs5jtV52RI10FURYfGQeaK8Oc7LGYsIXLEBIHacJr4sQiArq/vnVwrFhK7GZe
KCtAQ+/zJ22vtleL3wPGrYn4ADSBUf6TcZz9VYPVaBKU0cg8+w15jRP4Ic1srLkAODBCxewE0UsQ
TT94S1+FERy5FgtPotBE71UZ6MMQl6RNbYHKWBZc7iGRAAyA+jBy1e21MF+YAIrdCF6kORigq2z1
Po7vJRIS3ArFmzw+8y6EtAdMRtcukNcikW3BZ9Z+l9qFza07Ndjez4ViWxP0g02rqdfcB1hVeVw/
bMVPxp/JEwJQejBGvmK8As1TBPTtBN2uks9tcrw6g9u95bkRlHqWMK6SsOT0k/NX3O8ds97rjRjd
GoaHEvrpbWYPaYeNkWwTEJ6G0EZtBgOqP2LogbvvCrx3bK6zdkZvajGzWbf7mnNO8qbqbzaDdXc3
Pz9JWXeXoK+yEdDeO/pfbSLWkF98zvPrzClM6X/Tufz+/qIw8y7DLvpSy+oOnf13772wl1leicne
fWKPWrRuH4J1ICybCmHlb1+dwnH4QxvjT8kNjYpGqjn6nAjqsMReptX0gtZPBsuJ/4pjRMAF5YO7
9sdnTsTBNk0tjfOH8xRWFn7sCFOwgjIXoxPgz7okNtEcHPP1vstV9lWWvFaH5E87DOW5zjciy/Ny
8Rs87huKKkyJ0O3DxHEBy5vI8Tyz8RzJQ2+dT4rzTfVfB2xvWQXhxiERjVOmkNeiI+JCd5C3RVJB
qbYpCdWlyMjS3WJayi+zWMD+3BzhyyVlpRhZnfu84XcbiSiS6gMPttz6trfTH+oH1NrMph8DC8dr
d0qTdes/u2Tpk/iOvq4/Kl9NUjLMWIzfa1beDdLDs9fklTZMekr8Dytykp7YQ8fnw3NW1aHs4vdq
l+ayRL3KjBV65divlOUiOGy4j16pOQJECtxQdwx5di0eKhSWcm5XUd6dPqR3V8Uqf9q2TOs0NbVL
u1U2nnMjoEUuClRSqU7gTOId1gs6IJ+i3QOaRu54bA5jIh1BwuN3wxrmMRDVQiPFKLJAdqRK/bUH
/YpBpb5UlrLExhKgJ/u989ig9CjTgaDqzcBjqPKRTn9GhnebXhbpL9At//iYIKtho/WHVv2xEQPP
bcZMIEZuO7YCfI7o+pIY8lG4qm0toR+Uu6Nnm8IrM03JgonCigCAzsNrClGGuqzQKwdDTxsyxFXT
yVaUo+N+rwXs/exK9/sh7JiKJZWjLjUtlfXETfJxaUrJxcCV5DqZV5Dby5bsIH9FvfGE4/S10ipU
e9Md2hVApQNi6e28cGe+T26enFgPFmi5z1sZRi67iVRMf7wa/oa+Ad87clMLlF/03U99sc7qDsTB
G/io1+yjET/BoXuAYZ6piGpG1gwsY5Sa51YGPFJX+u0P/iGSYmBcK9zswH7GKRAswFE+9/t0DCO0
gGYt3rz6LsZN0rBJv0747Vc3Uxnu4LnXX3bA0PnD11JCAVY8dSNkv1R37eTnakC4Y/wTayNMQkIB
InmVx8kAJds6BCDzkGdDb1Daxzx1uT5JmVXO0xb4FaIlNPIPicjDMb1bOsT0B2NMGKW7ECTMAkYK
sh9RSOV79x+1nT9SfvAvtbFrefvgGUuBSzGmhYPRFYZ2C9MiTFkI8Nevha0ZwsXE6OnQg+CwbccP
8zuk8ovGePr0JBYGV5owxnmSQAPN8pqujv2AujTrTBaAbWurN9FgY/S2Gp1iyjeT7rM1fyJXGHFl
FF51E5yTYEfp/CHP5PWmAPOGhzppynQUO7ftGPacRCzWzOT8WT/nIYHJXuFwH6utH7WqnLCtabS/
/YfM0YV429hGO6GYUr/hxonp8A2ArKEyOaegcB6JThnOVD9NOLzKPDuvRH0An9oLkUoTrfE9UqNI
MowdkKDxwOf6O+3swL0cjWtziqzaWm7qv4OcGL0OXS1KO8B9lQN6ReM9CZNrMODw0zl6xE/mYDr6
seX3631Xdpcjnm0GimIy6NKcCNozPpX8KsG+fTgvXk8XYwK+LIokYjJ4iiNY66dGSar/kgsQ7A0o
0T0SKHxmvjnN9Hxjyj+aeBHUBsDwE08woXaDCUjE3UNWwpe8PRdJi+gkX0Sw6e9P0SULtEAHal14
/d6xo0geA4BIjw4R2vB4+di7tdeEPH/8n+OO7o2/oog7jZbrr8+49mnZL6ZEd9XoJzPO0jL+M/eM
iOaXDzdOfTFkLI9nH159sRZbH7Hp4LB88MVdSesRDVsiPp843++nLbHvjpMDUk9DsLaVC2YNaqaP
D80IAMHGNKEdLknNyZF2mWRrQC1F2qDvwgz2M56IbOEQ7ruR8GKMFKyTSMBm53p8g7kOR0oXtJcI
pg7lIPWviJrsf/GO5xt00EZCHXmDkDVI2N2GPtg++BHGUv7oGpq1iLTUjENx8nojL+XgLTSEN3Uk
prqEBNJjzruND96kFDhNHTGysve+CLM3Ug5YRMREAOCTd6PcURNdM4Pzq479N8zZdZG6LWguFrpU
DlZRXEKcazjshUgmr8+iRz0QwSoMgwEdd81EgUaJwzC/+VwQI574mdR0tcdGWmods+LvlH3wEEyU
rGyJW0pVjXoYb54EQ96yTDR+wCbIVARaTOrb1kJh770cuSamRFyqWSZNr3rzLLSEFQTZxTaZ6Xaj
7oB+fFpNJohOhmk64OEbPgg2UjeAZmevck+z4peuPjtffMTg+4XeZkdFTiEx/8l0eUvUHdKmj75X
T5r7hSTGw5fk0Zxmcf2SiN4Lt/cBTb7yegzTjt7eYygzcAdaTO3j4L7DQI7e3XW+S2toY+lf5MYr
HLWHuI0LHJuc2ppiKjsOpyDIu7ctqWs3bUdzAWU/xMaffR1PFu7+1a6z7Sm6jxAWKQHdje+ngd7T
E41reyTmyx9U5SK8PFxIH0YxrHk/oWvej6nrS9Z0hVWaPikfZbTtQ0Ul6y8nB3jDZ1xX9kq0Yh9v
gMhdzGUQw4YIPSq6LPgHXNqBhy2rh3I8ojdlsHaITpyef9c9V159Sl2ZVW4YKnWtcGs1+pD3NV6q
zazNG/fTJpo5LYOPypxwcgtetOVdQqLgkfOVAZS12DCS6Fnhhg3JfYQcxrXvoUI9CHkU1NH4uMFb
Hi4IpGaG63WRtOd073BZNniDRpbfNIVbOcwQSbgQpkjE9IMthY39DS0c+k3gPEHxh0TVYCZoe+0H
A9urRY3hEi0sQcFBgkcbD1GnPWIMmGV7MvirH3YlV+Jay+33i+b0v4TjpYBhkKsz96+aVqTMg8S5
xWvvmm4IXyqy7HGsXIJLii3JkyOsdJQ4Y5Nd/Pxbg2B2qR6W1kNLfHy8arm8Rk17WZT57c1metDW
NIODYhxI58qiBYKCI2Wl9XHyoCqUveTJUC2q6wu24PKO+NKUibNTtL0xCHvhsxKimZdVud0RYTmJ
mczAFtUGfkZuVZRZ7mYgbHBnLPqHWY5k0LobpLeQ7dY7JYlheyEaM6gQGqnzj4Sc7Q1L5VB2sUpZ
akkjF18kAcRnDHZbAJDI8q0LEhMJ575/9Sq6iQqocDLARJXJGL//+8ZE2QtJT8WfFwHouzdInPoc
9x8ApAu4F5RnSbqsI7QTOgX5QNimVxqNi0LPHfOernjwR3Ees886vU9PmOhT/iC2aT+0FjoVM8aJ
MR0dy82nTjcetn2NMU/scv+yUptZGfQW/cmA9dx183tZC5sNyeenKQbazjxi3A1PVXIfZgy5rbvQ
FagBMo/c11DfMUwQU0h/c9p0Zx1acRT80Ewmy5nYXapfju8GVWUkNdYddv8JMLqtLmMzUXFZHnjT
TYYwLEpbO56Q8h5/mzhRDUFFTRVbt7yE11I1y6DM68NcApzXWAZpBvaZfr1nOahbFy+ZKJMq/Y2p
CW0D1CT9B1lHv+NBkascRr6D0DYrEd/6BTBB1/Sh9doAxTeXsKzrutFWR7ANYBCLj5Tidmh4fpA1
NNHvbkcyksBtYpj4hU1zx15FtljiAtLpcNGD4Xxb5tIX7HsFmc9KCbVQmtErqgkItOByLOUAl1wj
QUs1KF0P2cUspzlg1Uez6cpVb4bpSy56OzF3kJb5BHFCmNq1xiOlI4Gr+n1nCdJAd4744GuA38V3
ZcG9N/zKJnRH+LGHzBKjpS4lRmkJV10dsP1ImNPGECeGQxv7psbUsVvQOhdRwImaggDTZ2HsjlQJ
yhFQxoZUvNz4CHveuNQ8rIN8Mp4v8NA9X9lKz1eqVceAW8KaFkQ4XNp3Z347tQZVTqE3W5tinGY8
CoU0JFdxouRZ/I2/UZ9CuD1sFYLBQFRx5SlBvbL7lPb1K9EkXFmM4ao/M580zNo24mOmMjIXUR0J
dUAyKMtWmRZV5bRF6WmVUF/GeJL9qtR9lHyiN4qx/PJj+vwOgbWNpaBtas0pxHVYaCI49VNss2b/
1174tAXpMYFPTOchUjSvoZ3GhYOLbfSmEI+9uSSG16+JKHgQnGwmPSZ6SYzGGPBcp0Dih8j+83IY
60Nev3xE6/5CLpbQuNSdlPRcNINm39xRYHF52HatZKZzKnVqQUGbMLVXTSJ8j9yhWkS0tpQ4T8tE
XtTycujcfkZ5kWbXOSvVB39NVi1pEnIGG1CX5A/oBTrQ8jzTKgaFw+/TWo4dMZmTtgffX9wjqpgC
uK3da+XbDezdaRcXsF2a+4N3eXp/BgG6S3fa6vOiCpPMrDCTQSd02dDvrOxYwnjKcuemFDvvvGSs
kRRVUez+F38Wzn4s5TLCvXFs+qjPAORq0HX3MAPNf0xhLYa6LfhLjPcxDFlMKG4Xo9xrGeYuhrdE
tuk1AiaEXX1rFyGVi7XEeeP2Al60BtHCw5u8cMGtauTCY2ZNVTAOszRrQI6YEgghrRNA+sfDjkum
uBGCemQTTSp+p4xBUc0ETVLdKmuhatY0ZwpLIAvzq3i5OZ3gcg9Lpt4Z5weH8RSixnkwkCvHMvFD
tqGtEOV45NBPQFt0RkQOrdaMhgJatmc8UlGWdjlmOlz8QhcL4RqOWmB3z0tEiCKMGFpM9DgJZ5ra
y/qp8vrDv8A3sY+r0X0w61Vfwf5Dm931W6CVgXL2D/NbMNvhuCLKbuu9ltGEEIWcIK/d6oyg2lK6
zWhaOlJvsjurBmRGiUZYcoi+0Y+TsGluLcPRlxRPA7HUkoiKLna3PT74aTWP11esrI6usPav0j8R
CUZsFqcoeMzibk3KrVk8fiPgDNoAZM/9CrVz/nqd+2lzTCS1hsh4Z1CMxEd5tGT6BVRmIbWs9c/5
eZNyq16D+g2+aNz6GYhCoTaBi2uCPdcQuj44Y5zpEy5U2xRSuTUZZ2BqHsLyQg/LJAgEJFRD8lod
v/LcU4KruleBhH6XjcxQBXZjSlg9wiuua5K/nCv3uv0CYHa25L0ghzuB4vvaylWJaETIhyDeQH8R
nRtDc+mfKfE+GnQ9HBN1AOTs5jBwH2W0mF4i7p1g0UFq3tI+dwO8tbmHUQE//wGN27FcXicka869
ZQLTAMfSdrYXOqRlnSn81YJ/pIlomKHX1APvBp7Lh+V6Z41dVIA0sczOcXRQvbC/xhtaGyJsd529
VdnMi1ZjFyACFxBJNqvfvSKRQvGtvY62XkQP4LdEN495eiB9UYtw0WonBawzOTxqzgBDcpEEtqVC
2IYd2RwibeK2XhXNoXWkBnJ2C6Vp6U2rTx5ik2yH1y2VlmqY7SMNQUPJsPgQsS6SlSYOT1H8+PRX
XOSdcXCSHAB3r7lNpPNVb3K7ioYfH3f5pTwP5fatu65HfusiLT7KQ7EZ9lJJsiOx353p4VlM04Z5
0KhmBi1xNSPzxW4WScJjhO9Gr1gz9MS2YjQT2HRnEvSDqVn/R43VlF+HhQmpJqxf3XQrLDhuUGIO
PNxJy42JVptIQug15dVbYFmJwXv/wC04Wx58Q0ViU96/OL5monCi5PpqJ9Bfb5ibV+0XqkOVi+FX
ZglYowx0QpUQrBUYoUR9AHe02YO2DxlXjC86bsdt8CxeWRsakn9B//q9WUPg8AC1QbGr8oS0h5kI
qslE5KiC1TgQvf5bgDVqEcuSvf2k1aZxt+kRH5DKp2RfKPFz6Jk+XAZ6GJ6xRNAUmUPUOGhioQNq
QMAYXUtw5nR9RlMnolKJYd9Z2qwm6hWdEheoY1oovUv6qOflmiikobSbE4dVm2TrB+capuSBbwE1
pmL4l1v+fUW3RyjA0QotRDRjHbm7GHurvmsBVs2hFONParuqSWYKms+SzPAAScywsz/3j6CcH8xt
Dil6g8G/yImVX55P0MQgGeWM1BCGi5VM0CCsAeLM783TMeppvL68qqbhqbAFjBu2NWwB0mTPJbyD
cEuGYxQpbLRwsrlu00We6UUyMjShLevBoeJUSIHRqSsVt9amtiE4rgwZXMLjJWUoJr0DFjPW+dT3
zYTuvl//ekUA+XQBuKSd6lahCe+HrmvdeFEN33j0VbGy7db6Z4Ky1ahbExkNnurx5tjCVL/IXtRm
QsXyUSgwoQS1YMSrVpDKCQY7ZNhnwNH6cw7emkdl1VaG2O77mOxAzI8feSeNwPolLHWqy7kRd1KO
HtEyU2FyV43McXsIPoyn0hwwj7Dopz1cbZQgSG7MyWh7RpBi+2Pg4miqVPagMajJS+W7C16nZpZL
wx4e/Y/3KDM4gLg2a69gQCRJCTS21NH4DmcptID87vee/RfhGH9PIpbs/Q9pv/sC/D/aTSEMZKh+
wxtBn3zOVQei7MJEEpxpaJhgZ+Wbfp+GayfUcojdnha4WLnYnTziXVFXiZQOY6Bokc17/2cbMAd9
PgXfKsV2Arktz1Uf9pcNpHbQhkyWCiohsXznrwBbAWwNP9olH1wjsBjI9YTjtdg+9MSX9WbQPL7+
/yHnyGghcN2U/HpXL3UKsf7ElleUkEhkYHBYuurIaIeaSiF6Lhs6YPXjm/fpisDRzghhuP19KYgI
RDKsYsu6akfWAUIJN0plmhetnLaEfpG4nJYivxqouhe8+v49g9acrKD0Ab15DENH9PefLUfbOxT/
WZubUph0yP6d+WwG1y2BVFaqYDGiy5Na5SVOQiAvJku87Boaqe1v+smeYGTIx01J/4elVM+0mvnF
DcdvEBtdEzpc89hU/GRIbwAJ/nJp6kDLkH5m3eeOuZAr4OcuhRVmLUS1A+tMc8hgMMRzLWiyrPW3
te2q5eFaUpMYKEcAQcG4gGhnv9tBKrBEq+8DiT6WL2EOHhXfZd1ZRjCobYzILO4ipxRJk4MyjwIs
MzZrl8rOH1DQZGHnUGx5P/wfESUzNXmuxHRGKHye2VUdJOKJ7hQJ2vfJ2dbezcLSxUlBPAinltNw
MKjqzkr4aAiRCrq5DZoDk7e9AcQjr8BvWCr46HYCljP53IKX+YAd7zZncmEyyxhtbeWAeIjxJN34
VctqpiQMol2LiwblX7ho4x+IXQAwmYfcvW5Rn6hq+Uk66VcZb4FYcQuuorRwFJi9eo0F3V8h6yFK
bTqvUajbDb3G8kdwWj2UJIy1B3KsuQiFWAhj4wdJAfywpLuzpO/G+ZpqgnjIFW8UISRvOw2jB0AH
9G5Ljpte//TbIYzj/brXDrDXnniAtyTvduQmEUTE7dP7qKMgdEBoSUnKp8xGQYKoyrZxw4gbawOY
b2B6fvTV1bExrcXvVW9Zx92qsstbSMO+smtX1XQqLfMaiT8sIYwkCvb+R1j7CtNjYtBth/nXkgBv
wODWQ+JJuiG/lzTqkPP7tHGcTkQJcO7AjqI9UbDHNlVkPhcZ1E7vAl+7hEq+H4noNZo/ngGCVOfg
Pa5zzyd2a51l1gPItZexa4KHjOtq7SDgeAiAcIjFil5m60JmJ+2qZqHL3ahG+ygPXTMyfPRoY8zK
uGq9k3hAMFAX9dnJrUu83FEJcaJaMVVmY6Uj9BMPzKEC+8efrloRyLbRZOOOBpS8f4IFqNOBzGOy
xEYZTeI02MuG6zkd0lGPfyOdo4kT+xG0MxjtL45HPzgn384VU84evD8yfFF8R1iiMKrjyOuzxt/+
zOlvRdA2Hh0fGqtOf+4eWQGp9LT4B5lvvtUL5jaZRIpJbHmfBcNp5FU4tXRXYl9lCDf4K24vp4XH
UR52Oh67G9WzOE2+7DLNIK6vIfmgX/dptJ7+6Hgf2wY/9PnZ/JQJm7cBYR5myg079tTJbJtNIrBo
oswuopdOqtvkYai1ZvMHvoLHVeI3+o4gwYoPFbyDSl2IHsxOdLQD25vqsNG+MGH2TfeEaM9LyfnA
wPi3o61Qv8RoUDTNfPEM7Wz/9/ke3798/jOENEXj0pC/152V3zAlKw7VE6FCW+TY0doyvW6sMy2X
s3W050c4S9f0n5Am7Bcp+ithQ3DjJBn8GPo8RqWxntcJkGxlUWawKpBIs5Iro6jmHRVj8W1knIJo
Iop7L79fEisj8V8ferDSjXLRBKRfIqP14g2FVxDX1KyBooWzdvnk2wWi38VatXJPKaGnnmsxdX9q
zyLRWkJaa0scfDFVccpD1tjNQ8H9qGkAH2L0ErHGpkkMTHLU+D3dKrDRP4AFkJth2HIcihLmWVvG
h2oCW48tvDfnvNEk4wyC4YWeRJ6trH2fcy9JOqCKyTjmzlDUYO/nxh4eRLt83qXYDvnQTFMGVP8I
B0Ezhv0BI8ZiY5JZhHiCZo2Navb1HvyBjmYdJ/MbTZsbUUl7BDrS591USbkk9oj5HkQmKN+jomHp
WV5EgDRQBFMZvKtO+gUltaaWpeVjXEZECM7T8eg2nn659o++8VdV43x1ZMmAd4uPx/SHOVE56eYg
7Ve0vtGymsKPCUXSMVzLtuEkAamMklZDIOGg2AsiFd9Heb0IY/VyZoU1qoa/5IklC+8lzQ+WKaBF
UE0IIRaCIMq/N9po+wW2RbQy+IwIafYkXAbB46gNkGGPOi5eL7+jWudeprSh8F1kPTFUqhOkyrV9
Ab7bGkwD/HkWO/9/PPQ8sIlkkpaTitx51lPAriuuffmDdzod0wwMfIYWkCklLgbdlTHQ/ZM3Frzf
GziZh+3Xgh0gLITvPqXtbDxAydyCMVJzeNUdkLLfQRpa/u3Sx+mpPokAsPuVmIKEFFsEM4rNXbjF
FG2PKzEa4rsJOQb7P9Nv9v/FGeQoI61mBQhkCnA6EhIrPYfzYNuQAgY0x3IrUJqUXOV3LaGsaseE
oDC80nlJvXHZ4Ljh/dZABRtq0Tk004pHtS3yF262N/iImDbjzrmhdGzBzLP2+m+MWkXhq0fUnQuu
QTgCNEmHW3dRnNEHr7G7QxRTiI9tjhGaRUMBHw8UXAZam5+Shm37QCZMjau3Gv+fxaSLDpphzB/T
jnQlIblnMyAOP1fXmHh4H6DxP78PZ9K6nmVD2rzr8V8tnA8TQl/E3mg09kFeinXgf/HCbNw2Rhcy
1WldANMsT73w/WYmHQ0zKqjeiQfHbJd9dNCBYxFDAkKsrACxr7c+K7tTowZxiSB5grGORFtV6Hxg
mG9G2I1Ie+7G0NEpPEc8HQxAdhm/3mPCPG5bXnad7bqqzVMRnm13CLJQZbBWbi9f0/5n6HLF6nTk
byP2KhkSx2T2+SY76CdpfFDWc/0SMVdL/I/A9M2DegVzFZo7i9zh12GYYywlzNXZnUDMwJIoQGb+
O1Pcsw2Fv6arIr+q6Fbwr74Xpc3lBpeOa+7EcrlB81Kqv2eodIuxO+RU/Rt/OyEGmSwpaAH6WcSx
iJJ/LbZkpJXpPkOyJdHcsdnQ/0jk1p1W+sq/kwyOfeh/iQwoHrhuAug8aogajIx8vd0SoF2TGOq+
pokoYcNzM/lg1bX3vc71BPafDrNpDNUxoT/oCVQCxZgODMxtXZ/qpyF2mv2Yr/DV4JhFsDpT6xJc
lrfFNNNW1q6+OO8dqJ+N7GiQ9pr2MDeaXFEuDBZgEvWT0cUGUtYtDu9klrZi//ddUgA4liZepgD/
mF4aUnVaWM+18r2+llOpizsHVhQhC2mwvrfW/E3p17PiBbZi6QDGdVayMXgeqfFZZPKYEojhc/JL
4o+ynHbCKrWtn+kurODWZogpjBx9pOyN6rXyyDzaVfXF1t40+RO1VvLzqJF/SDHEh8FDwqXIZLLN
FiRiKNRVlj1cRpQtA4SYZrJ6VWVjN+mxEeYjNtDGm8ySczcCnXRt1jSmoecdDLWqbwHMx3LC0MCc
PDoBdxP5jdzfx25Phbo8m0lKMa+he23RG+5BWImkFIReyFWJwWedS9WrHkrOJpuDXrIKtqm6ggx2
f09KJCkeAgcuzKVfmOL3ycISXQos5TkBXNXyGxKAsihs3cx8EnXg7hWr6x5WQvwQtsEK1Yq+vm1x
oaRdc7ebp6y/hYIml2Pei5Je1LezGmt4NJN8aWhDXqFcCErxaje0UfXiqJ/grfhMogjDKsjXPGsY
YdE78dx+2cv6CqhrUOIJy1fJseEQbLyT9CT3hNTJ3xgpSdCYV1sas+zZG/nD/Jet7ApiUSj30kzt
Kcqn9AUmsgXsgAgUgoaOdv48+zMH/oLAF7h7zBH8u0u0bb8xQoZiNO7svdGG7LNJNi1M0odJShBQ
+Nhuyht96ITIlSu3lcICUGisGHG3SSYNJodO8pdwcU2gpxdikJppYsk+UKbT+Nu1SV2XDWpReBh6
iG0Wo+7HZ/lRjp+iGj4Kt59y0ERSQflXQqUWYl7beC+LF3Ueei8eBR2rN3XZDC2voJgP/Sgryvh5
tlAtmOAEjQLaxu6dr/oGDR9wf2ICo5piR3LdvZN7eqeiC9ZbZ39ux8CnIEXoTWD5/Lj4HpxDK1Rw
8klUh9TgJl9I0XhLT0Cpqguzyk0J0ouQl5u04Bd04vzn/LBC+i9VY0+aH5Q4pOT8CE2gXbMZqfd5
ZqwoqczIOrdj4HX/FdA7+5TtgCPxUjcpet8+PgMzPkonYNP+Uvb3SHSYKony7ebegGdWFfC3T/iD
FQy/F/ECNeEb4oF5hekYjUvK5KRcT3xtjjlHbLzK6OtOEjdeGfiXC89DZMUWMHsJfOwLb8ei/rTa
ZWUdujcxgjc25GQJbakvUg3P5cemssVRpSLEu/QIc2tzPZE771H2AtWq6IE4q7stY21xNF9IcGbY
m4vFGm9hOLmzVXqw9Ik1uboWWLus1Lj+248OpzC2Ji4fWCdhYxanua87J/yrTfo5Mj7BNZYaFrHX
XfKvpkRWGp7XUUYwwUQ7Bf27FmGaU/wmsKxvSEuUiXvv1pRIySRDdhceHn/H9H3YyssSRGdMSI5q
vpallcqIfaDhKMyVL8wJVdGC2Xj9kb3T14sK1Rdb/lY9Q+4hKU+pDLUd6oo1/KoiU9r8/fzsSig1
NDRBdEHtjec7BxWBgXtzB4es4gMohsCaMIt5YJU+qP8xO4dHLUnnneBd9BpBrlgKzZdcsZieVF+H
MOd4nMvVKmQRKlt+8u4jzD9NVLiCB55B4vNflHMvItABttF9QZ+pEu0tuF0aNKvoG8pQaKTBcK5t
E2iK0MPAURH1tYIkJtS1xnRW8r4PV9XCYQsmUjbWYmyo661mW/selcLgh1GY6fHml3QvysSLMBj1
7ybYV7NMKu4RtY0vuqmApMHktakOouMW5KFu1cpdsP1O8gEpoCUTxpnGh6ki28UPFS9Rj3yJAjRO
g1rR25MXF5TNFa7xtygGD4Q1+xWzugeBYBcj7CCUd3eRXeTql3aE//MY8JAEV78aCvMDYXllRTYS
vAnKFaC6Yt2SGnfUrNUb6U8kvAMU74+c+NWmR3q7gE2HBMBzKKbiVZAHzFxS+m2g91u6Sg6mXy+0
bwYG0UNWSpU53pP1psYYWD2WffdVSnA8dpYFEp+BRY1foU/YkkIY7yUaY1FEQRH4J76lZpQnY1gB
eap5gzaKzQhnaDaXxi61xMZw0wYQ306LbyZ8dGm3NZh48TZjXrGEsiV+CgBh9ODThPfCLsT9g2ju
bczYhiGxM81uAP9iozpOB+IvSJjM8A5PZMhCNjUNVe8mw8zylceSWF/TSL9R25VRcwBoI6KvSIKr
f49nxZ2XbO7dBfPUfQ0mJ5p4iUHtRFvkUW/OcsbFmZDw0q0FXDnWNhiRsxoCDvuA9eGw/uEGxXtX
3z+F7tk/bVTE1IO7saFWAkiQ6sHIGYLwbuG/qbOPW63ttre+/JOs79eMOWDfyOEquKEuBW6wuiDn
U8Xqeg+cfgVD90HcTbLQPhEKzqvrDUjno5mT2JHTDlzJC73LKmAx5mqmDLhgIeZLrD3RIiEBs9BF
5R33MG0taJUqEvy/DG8fTAXYiYNQT74w7TlX6jpfvVwW0LO982dgiDDt55TR3moy3R6Jmlt8QVxT
FxMLnJn8S5ym0H7ndXSjX8ZTO8VSX9G0dKFgu+gB49Xb9uCO/228S0cThxW2ygChiyi6VxGDz01H
UFoqE6+yHea5KWaRwyGgfxZnBsBps4llPlVT9OI6JGKXcxyKfFe46F3HigKpZrKds2AE8vnlfsDw
3WRcCPiubt1foFyJq7urqnWR3zjaOJJVdCSW207GXptfWWEIKBgUybK0ZYjZiHzZhXce+IY6j1n9
bpdrFX6XBAaT0hQ2Ntu5QpF5haZ4mLNI7RMLxPDzWE5qCl3F481luNewTFmeai7+cWyI9T8jGOvL
TshxyyBLee5cTn79aAJ4wp03Z5KqfjDAZzCOkxyNNLQZ7VFzFDWf7RrCJY6Q0xqn3i/6pIUOCMod
2d4DcSAcJEj5tiWlEWASxd55yK3BSmxHWOUx5Gjd5N8Bphe/zY6hxJ817nMgKoOc0+lknDYa4bvs
LqCdN9EQQDeertajXFNL3V9r75FZalhyXzUGSDnaF1sOZLTaSv25OT/pcDV3fRm3LH95NW3hZl27
PPgZlMB9mwMmq8vu4gfkxyleoTfj/VQHRZm6HUPnBcpG6pnhwNfaEHeLFAiO0tmZGBrIrXqve2HR
wO8uEfsVyNZ7zFpDeH0E02N2wugwJsGtNcLTavkChjJKjRFMEIpsoMObgcdmg7pLscagyl8Uo8ND
LQU8zjpLRvzbxirZzmx246daWbHq1EPZKhaKKD6W0haRqDz2YjRslnY6UsVLBPzcxnt+M1a82L64
sou4Dlmuc1CpUqi8PvWQHM96DL4Azg8iHPLzJr/MRL2gzwd8OSqWRvTUHgGbjkn9PTsqcC+t+YDG
95VLKGdKlhYbaw/e5ux6I7Pat92n//Pup4cFhcmBasgb//PofL1AE88+9bN+ZaR4s2Z0LJzDYkLq
RPFJvguzgk9Ns/QMc5MPoLwju/F/r2LWDJRB+S6Y+XRBYLPnpVhOk6jcHsW0nsuWnK0kME3d8lVl
2SI4pQkCVSK1KKHnzZG7OJ/vw8VjaEghg/70rNvMG2Y6aUUYPUdFH+MzXezDYuNGKWmm0V0QggRN
EajVLAdQBw+d1DQdkfWncpxA8KPNjABQFRlRW1116emUWhT5CY/NziqYXQU4IaoR9R4vQd8gudrF
4qwbwJYAL+Xht6usziVG1SFZMU+p8zlcYs3SseU6ZXiA0EdSrUceNmylSQQXWmg5NYRjSSbmGn6S
qryP4Mw42YGQkGgYrTR3PNlALccAlpuRnyEo2Kv7qYAbzALhy97W9S3PkKwSvOI5bS0cBQuV1zRe
ZOO4BWxqhd0cN40qi6ixrGVEI9VBk2DvsznFYouVgwgy00R2SpZKhVmQdEBjTT7UiXV9lh8SyCSK
hegyBiu+g5JIrLM+fSGWSvf7qQNNYwBpBoOv47mT+AzgsxAcRUwE+iNl8gi7zrbMoi6IvPGkl6bg
UgGzvPD/xEhQx3YEEkaNDLRYmXaWkZyJwzcSN9p5n6rK45X/LvXHivRKTQNNREboeviZ2fp7pyxR
sJB0H8S7ZSbv4cruRqdI33Ft6GwFUzEwWmmP9LSUlXpg47rZjrUBraT/yTMn4EdOFwj9MzuhBgi5
q0NE9A8nJGgQVUdmA4y10WV3pJsWXfaNsTRBZkRvgzvrb2BdtXuU/B3KLSYFZG7MB3lM0HVI4vXO
j9oYbVx1vaESr2/nGNPiWuw8nZ9KCs4/6IQG3EiQiSZ0EL0VEVH44TAHU0yFB84UElCAcHqkhzhe
olIPMsdRSdSKmfDW3OqMFlx24S/FadNmWLBq15I64sU0pX2zGQpM5W2XQPysZ7dlRR4Ndgbvi2y7
pptyBGa4RevHSZ3GbUX4zHY4OOpLWvjZ9ublweDzdZ9jVcWwbKh6k1xewUnzSocceC5mrSqHDOTk
TqFVewQycr/Gv1oZGmR8a2yKtO4w9me0e5mPQGABGPl9u+bAYONJhOXeagh2yDF/n3mGk8mnZA0L
tx20bb3PuqdoXvmZpWoHiZ/yoUCQQLdAsKwYC/UNx+UK5NwsO62qKOpTRUf+zI0mwA/yHbjISUXz
/ogLsVdTLrKuFvy1vuHlrSayf/GuX5n1+4881z22m8ZixcmQsFA2dqPtukUgh8dxIpkS64vi/jCZ
alFWQFzCdhlcAsWSmUWn4QAlbMfnX6zMsD2Qh6LP8B4E5XWLK1pVTv5ixM/Fo530p//TxDONfX5L
4qyVf5fEKtuJbhDVL3ELwAr1ETw6LErQ3rvBDiDIZ1alqVA6e+PMa+YXlp6a1q3kV1dVaJ0h6riL
hnp6FveL3uufNMOa3gLIpgzZTHwS+v2v99dNjsbgsEFfmtUkPW8tCchbC5Nx1lXLQjAMnwGQXOdE
tT4Q6GAhHKk8gUxKWwcqYJKYvPVykyZvXU6UILepMcPqQS4su1AxtYcliDthmfhOauoSVkxv4Kdk
WmssnmktwFUxSl1kGQVayiegXz5t0OqEmuq1TDpwtXIjCID3PQHw8Sw6QDjP7Oho+fT9Yi+aF6n3
7R0bR4gX2e2hKNJmHYCGPcXi5fNV9TDjrF5C5FvcDKjQ3WA14zZLrBHSax37PiimAD1CLZrxqtoK
uKCOY2T2FTvE80KL8xqmtJnQGX2C/Vi1euUKI+/S9rBt9Axoclg3pKqGrrjAzeLXPvNu8Px2PTRt
lMhuSzh0F1lN13AnF0q8FrQy7xqN2OZxw0jaKdpTDKWgFd945v7y7RqxszfuAICibsyZbz8AvWlP
EpDfTZZ18D1gJj/ZWswfZUqZhUYi+uGmrX/GDPpztOfY2t6GELd4EAwqKvelK/mX4bvh4AABpu9s
V+6JejSA5TmvV4KLp8A3vmEz38n8R7Hnd3slawDUYDprKgZYIGpNitHSNLp5Zh102sdWahP9cXry
sFnDJgJiDPGeKjEJLFzjwcvXLlTsJRPVNjNjw0WOHFDZKm6pfTLSVhV/EXCz0Q9goEb5Se2Vqo3F
zqv905aIQE2PkmQ36jUs8dRKbRypUiZ6uMuAxUCq6H2bdcjlYJpY0rvYq9iBZmASvF3Ib4CfXKWj
G9u1BALZO/LqXftNGWvqzvABtB6AYVRbNH1QqR8nkMik63KKZ0Yszv7WH7752hGJM9705+aqvLDn
aP/Jtc/FFcrnmhLnwiZkVt0XmFjbc2Lpe7G6/mmDMhuWZ8bCk202qLHLpzlB5GHIP20u/UoVGmKG
PjoOHv73XaE/a8pULT13835KTV00W2wV6iDAT32TD0u6xO2ezqwGzae1wLKTMhheaTi1SpsvivQQ
OCIkYQQRBTnCHTQwdlkK+9n47l0zQ4cxBIngn6f6ta+0dX9gaf5/amaRqssJzW99KFYyURczTNu7
302wI6Z7YJwFAmkeOd03XFYEgFkYSV2afHTsbixTwyVd7f5MCjfauCps+OrYlCUqte1igQ/QgunB
Tu8ZOK+QQ5Fa1qb+g0BKG7CpjoAfBuCQIblPQHWqUA+LRJB7/vXBfFgA6FfSZRVJiuZAte3RAn2r
r9uJUL5YKCtMTnClM4h0x3L/AfkwKHJMRB7VciAnRe7bB/jKrhpEgAtNx+n+TMmki3Dg9ECCD7jm
4vzgFSC3InGjF2wL4wB4fVRD9uaUiGx0hHbg+f6KbadWrvMUBl4SudtcTfBYIKvfy7LkfB5yMCKd
JPn/HdoJkzL4vgDVD8Fe20gQ/P81b8eKO2PMeo3EK7EohbrQPbkEAmmoe2wj250/zrEo56zMvp83
XWXAUjVDau02drBpDkA2WsyltRoM1bXvKDkbKYkRuV1XdTV4nT2GvMzUbFJ9z1EE1jYdv8deSwfB
yQKrfEQV/op4PHXz3xfiNL42enkr+4fTcxShImSke7ivTKg9QTNn52tPkYbKu5A6QyXlcjC+iOSD
dUlML/6LTEtGHz6wsbou9OYnmCMcLctV+UQsrvN7P3CpnwCTApt/nv7XHPHoJPeN1oFTbF3GvS34
WERLRfQ3HxEbeVVCJGqNs9JQ2G4bNkmgvTHO4BEjm4bxuFUKDi6qbuTQXW3bNjnMRRzkYD10xzBL
jFnN+PdOa5NciwnY3Bnb7Xk3J8HeZj9pzR4yQzAUMVTQ1xGnWgevuHLdoCeXmanZqHE4nrwp0cey
kl3TxEC9nFmI9Q4Aw8DcGN2///gWum87VMv42l9YtbJxK156vnRIi+TqJBBj9sLZzaqkAhIzdqH3
Q+QSRNZcnheX4L9Rx8UoX4Rr1XJNmUm9fjRN41567DgnZ2QBM8/ioVQv9XzzqdcgMUuV+kK2Y9V3
00CnpFroUEp59NQ4iVduM3a3Gwt8qC+AafrKO74cxqCjzEdRDua+CB0f5MP/YDMY8uTrnskSmXtI
LB2S+4T2ZLA/GGecDDqzWPu4zOBgrlSarHudXbQFGScVFUzf+xmVpnOYFejFZc8Gogp4PJmqSEnx
sdhG4g70FVWSjtcTQiqlJrR4QBC5OUIIzqP10LdqX85r+6fK7FeVW97aW//b6Gz4/ndUeXqg6m+9
yVEP6Yd5pdL1hsAqF6P2KhY7Tki+QPtzDFb+H13stBFrcbqHwK290RR5wSsA34QgiGq3kCM7KLA/
e7NSLFkfulE/fV1phSmsZlDtMX4ir1GJkTEjqtZhdTcIF0O3kOka64Ek5h4NIa6kqrl6JcRjUsyn
krkqoXzzLQppuGjzirphc6muJpJeWU0CHbqKMgZlPWIxN6qcYvt5uTQHPjIP2I1rN+9qjBM6xS/8
RG6bHwCMGBSwjX+qraKH0cMZuUOfzyfiT9U4vkgT/gciH8+AFuLbW9Ghg4Te789g8Dme7myAxENL
TrtlK6ru1QBB5tJm5W04QVyVNP3A/3khY1d/oIFodsXauu6cLmfDMl/dWT3XlDx4+9fplNynbSXe
02XP6jw+gpbV4Z9HRn+B0EOdtP0DOdV2bLRBJd5vFSnLXGKfqL6zWjmI9GkYruB1SxM7k6v2ad28
hr3eKNAbwNlWoGHX6nfWNHY1STvtR/BCC4zMJzfnU9dlVLGmf4+OXKmPoXKadWIsOxrM+Q0jNeVW
90bWQ4OmTy6L/3mT1CYilss63bKvFYZ0sJbRzJ7DzhiV7aMzKGapFiMbW/VPZa65IZCNs8h6YT49
UNu7atezc79qHglgckWfLfn+L7fHmlDqFi+ZMLHOJJEg2w1+Dhim/JPwtwr88XUKccTdU1WkUuHw
OBFK2wLWDTtEij3mAIrwJnXO4WOb0en/8sbJnN37249tCTs7q4vUmf0Fsm3EtC6VdeIOz5Qjk4Gx
0Pr7Q8cr8Y/Z5ZIUuM3wRW2xdJ0AM4GR0GNa0Ei6EB5hotXEiuqfL5dlMtjHMGmtAo4JZpHXc4SX
GcBkHS20bepQb/OD3m9SzOx97nQjZhLUeeEwYfp41EE2L5WGK4VsRvZuy4DeqsxJNQbhnwiVwayv
WDtmVw4w1I87VuO587NuTuVC7i/qrCGE6uSt86CY/bQM18x1LYm+Pk6sO99uNdqvnVXnZgLQ51pR
vA0KqRXZnJq8X/k38Qngfaef70i4SQLf9xdVLKTo82SKIpPTAUypyGu0tdFQsbbrhyu5zbloBIiw
5P05yK67xpMIWvXxcNqSGK/sWnePCKFR8Bx3Ept3zkustojnBXdr7sGMfBzYLtwTtrtPc14MpKPt
ipdKEp+Su3yX+IszMttXh3A+GX2Lu6Nvv20jM5Tn2tFh9Qq5fSychZMuTf6N+qDA3i7slX1Rfdhs
0a1qipUltbtg1PVOAl73JfXyZgfUX6rzuNduSl6iqSp6yOgVmxqJvI/THtw2f/T/imRVNN/ZabCr
wn9KPFQBLkTuk+JIwPbMEVHVPNi7JFCWS1uwRKXUxRrbLAgpHaMpt4ikKXS54nWcb7gkylewjvO3
HDI3YSZw7YECBdSdBUDUsVhQfg4hUxdM4nJoek9z2QOD0u7PKyJ7KnBcmZ3/fm8F1osjfdkVKmut
Jd4veqrGUquCfSQqnkYtCj9NBh8Rcf8e7aYnQHkNExbMh0MHBtwh0qBDPQmyb7Bod1pjrnsZR6On
RSTK9XbpyUhlzAtXdXlgdTK1QOtB/z1TaCmEv7BQChfqrTKmbFqAaGzFci6e0oV73H+/AcW/V58J
bV5jqKFNdMBhfFwziVCdL39s4jONZzceIdkRzr2SRQR5ly6coVclorAaEtm+AAsAkJGVHscthEbz
CPXnvVuCPGbBRpeQjRL+H1/kU+vWCMg0DlZTqgasvzbfV1Q+yiOxQZjr9HRFRZfW0CFvXOql/XFo
/h8zwHPcIby6BkRrxDsDJDpNnafkfa9nLts61SYw7cp3U5dqpXpbLyrVDrLHydSk60bFiKFcqrqy
j4oopaswXcG56AeIiCcldyvDRdolpc9H+6wnZyspQpIlRDaDjgQ/tvEtDVg4Wa7T9PWBIuSBu9v9
9mTUt5ZsB4Tu/xvvUDA79HpbemzCU2AxRP4HM24Sd+OHmwPzkDiOZXaBx+/EhauAjaCXmApZGcyp
TJA2HB+OchcNKufRlIKmB2SjIjwtncI6mLAIlRy9qx/Ts0WCcIVpvWRLBWB+jovuRKsPg/W8iQhc
Kl3QijAkCLOzJTz6x13IbAfKuvDndrxqHk9M0B10Use5Lv8hvnXgQixIwQp7FtKxTVk1sQuajkSv
PGCq3hkL5MfWsIoT7nvegcPA3gl1AN0+vf+t/IL9rqu4iwEffSOdXqTMKY17660Q6a5er9QCBRod
TLqtK9EUJbuAkOTg6pJVY/4TgQvGBtDk6GHYuTDBtHgbs0Zz1AcB23xDv3dEzdJ0vkI/iZNMmj/x
wtbn2Y7/IjF++q8TmXVxYueRmsvvMPVUJVmGmjhJDhct7gjEBCdtiVGndFh0g1i5rakupXIkTrs0
p4zJC5nOlZuM8pLE+QOWlie3GXf7WOkVwyEEdJFikXkxu8cWw1TNOVXjgYGDqO8S7WIofw619XPq
xbpsxCF7RYt9svND7s4bga0Mf40OmIfATu4s6+x+Rf5KKvMlyNzVipUsrSBHt6qLYiIeGaikqUJi
q7QZPv8ZVp1TH0zNY5VExl2KJLzRxDoP5t3cFp4TlegI/OQO3JFFjmVmor5+qpA20Lb3JBLmTgmI
+7UGB3lmAMdBqDzHvrzjbyBPvoqGNkykwpPi1JNPA5OPsgJP7yw5HxTN/vKaUzZUxIP7HhDAqzPP
Vee7I2OanoC/gSM5gtg+zF9ak/xAMDvMm/V/rNgUovWTvVMN0QLx0zY1XlyoSk4zy5gvPTnMoUix
sPW3p051pKFSOAgYrGjhJLANl+kSTEkMXtUPSPJyvB5GnIC5dX5VXZSYtquPIt7bIQzp7HjLogAv
HPCigJiiKReftqLrmgjG8W1lEr9HsZaivf5YfEEJABKFTShlJk9MqUl895PMToBEQQI82jytO2DL
dumsxFpLbh1t24sQKf3EQSGxM/3jz9wqtEblV7ygF3xne1SMx15xmELgDRiGY9rrwZMAvlLTkt7S
DZ5iluDvZGgOMYZXfVvymAeq6vei/3xbB0rRV9/iIagaCtTYXxQIYRA+mGW9wLRJUBSfzMCISK1N
EOfxG9digLQr9ANSgGPdXmPvmOnYZwWYl729A3/UPdBaArOK1H+waZg2nCpVgPNs+lap2g1ruDd1
sx7oWTT0BU+p7qY3Tg/93CjRox/f3X/HjDa4JKNmGqCzQ4RT1RB21ofKfQj58fHzAliveynN6H+Z
GMBQsOAhSuRrlJPL8dg9P7h8IVe+/3AEqD+5j8CFrw6A1IvJ2PN3BKaEBNoUwGyVvZfnu7UScbP4
G8M2Hoi7xdycBqVuVgcERHw63yWfyBiDUC6Ie2gwbltPLpMbxVJ/JqoEsRozgle3eMin7HEVE6UA
kd9BGyzkYrHuQQ5xCmMG5JXzKSFCcSRgqmLJduVIK9Ac5lyFcoxEQZP9oZAfRP17Olxa4lseOK9o
PhufHsFX3hZMFZ6gH07xxSTSQ8oma6ljyG3ymJiGS+sHzWEhOalok36tIqEMwBEuy3QFw6WUK294
fNJ2rtlhpyD6BClk46JZDqi29EiiSqfQuq0MLSjN10AaWr2MwPTgtW/zLHltvI0CYjQM6mcWPHvR
f5qTYSaxZRjrR/s73mYG8oSlwrWbShbTghsXAZakouVjsVfNWpR/ziWCCYN6zhFZKd40tVrEs3O6
Yslfa7egiaO3hA9WyfxyDjW/W6TZHWpQIQIBQ5xvtb+dsVGQo4M6E+IEO36rKi4vlOOYiZQBmBBf
qWBGVJgeE7nKNBpb8JPKlKLzqo/jbPYfoePzrbCNBa/dEMQSxpjwJQUaN4J6hWNwm2K2lFg4lTzS
ub4amtXuiBtwR4PU2pttndZ/nnxK8lJmZB8nr3dB9Tmjz4Ruhv/eHWlW/L4FvFBMCWVatY2U89+g
dZJl7XtFDt59MwT1IGox5Zfe0qEKtW0/z2jgcPnMOCQGhhNP1PNzJOr8Jc15hupwdoH2IfDm7gkQ
GXr9PMB+yasDe7V+OMnzPjhed9mDhT0M8GvsxhjwEIajnRFOpPr0+W2EuSa808HLT3GQtSSjMv8s
k7i7Mqzu9o/L+4y21Ax3ml/0lWDR4R7E4k/XhX0uA6LaT/ffEi/NQZdRQSaBV6aN9LMRJm97IF2W
C9QzyUWwoPKgVv+ls1AIM7yzeQ+oi5sy5wrCgDfCqj8i4El/C2bjReDw5tg/fCjmYVZpnXvUBAS8
qF5GMFGfh10AWqPnRMoN0uJIQUv8E53XtokQMryc1VECh0XVj4OKLiw9KRHu18cJ/F5vBDoHJqtm
IXFO16zwqRKJAEhb1VfiTWnK6ewkCRAQR7mYacc9kZH+zdSlr075ewKVcjpRfXgq14wWkq09RCku
QFrcNOKYXx1NI7x0tKZIb2MrMutKPbVIBTFmfGFSSVYuHc1vzFnYQdb33ULNeG1fWRjIYuMsS1t2
NRuvtC0A5m0UD2AFuqtDTD8MwpdB9+XUGTtmgqCNMydyZxL5AXZMnAiOE6i7HuC4ORdq2O2PNu0B
BNGjZSyDtwfdtqa78MbtUZs9dFdnbToBqknJFIpHo87nCrj2+0L01s2kppt99N5RIG/dzTF7/56c
zWCyyMOOriUNoN1Q1Rxn6zkMLADgesezaqaLM3bx7iZMgY5LKm660Q2Yohni6KcN5qNg9nSjCZw+
rOoaw/EGXAQ7Bvep0OGP9t7XKgR0v6a7hfuQ6TItSIChbNndg3wgZLRlw+IDFJydaxXLBXwyWkVf
/yXB5mMmZS6sBlhtVBz+KS9VBFMnP/Kl8Hl/S9TdWkSsjb8NkQBDaM1M0+IHAdT7MkVfKpx8hsEd
6E2fUv5Q6RUEX2rQpsq7r3lj7xVrVaN5IO5YBiqz8duJl4Rki1FN8vJSRmo59yG/YItFIuOck3SJ
IaN9EksP1/EyTxwazzhxTQqmfaOvZFrWN4CQG8tONDFor9uVJZrYfE6xaDEbT6xEKaMXvwPB5C4k
V+wRC0MVOSBCOWYElPFTuSoWgFG+CDOlkYZxInz/3VZzRMlp5RanCvbtO8PbbjM0X4vEEkIBNPj/
WmrZxYWzStMKxNNwLzV/tcB142TknubKSLxokcJL++VZua7ovKaN94hwpSjQk5bjIuoUgjnb5V1J
os/SObGczaXXUJ3z8lTelFtCeV2niIM1kgGMLuCp1jGsuvzQ5RFSXuTiUfgGL/e8z7SKTuk1YS1L
YTEsk88QQjQLxaONQo54Qqm/CLiN0WKjg5YknMpcfjcydDgmZ/fJqRRc3mWKHqwgU7V+S3Br5SDx
PhcAMGh9+LZ9jobaN0SErS6+g8VzgyY4UmGJum+DQ5dkM4Pmkv9EL0zFmM8+c9NhX8JvZ0a4laVp
MJvjGe+Ges4diGHHMGR4X9IRicEjK595NFuWQRJfztB/Uw7KJHK8kE2Ft0alkN03J1tje2VEmIsp
nxnRml//SI6RR9LUzWZJVojZDeWbab+zHSo+nb9XF42PmklG2H1GLend7cBekTj5vR/oolkir5Mc
Kg+tZxrxHG+NDKY+C5c79KDjWEdgqJJtzo8zsfY3adh/3ocSDx4zBjbh9QVKSdvk1tWk8s6fmRj3
JsrpiSfrtJss9m684QeJjZOEVR3moSDvruxqBU54LYbKaibPZeuBp413IOPCaLfyvEwYoE28X7UJ
0UUsm4/XLcWrn7XgywcYmjruj/Zjnd4Dm54U9jaOTK25uLtLLhQwS3KW8fU3ot0QOToVa8q+hGcY
YB1bzWfiluSXjuVKxkXiO9i/hJn6QYKb2aZpmZQsjSCSil4r9IPI4nCARTBNQy/f0eORh7qPFE9z
31jtlt1wKnzaplSk0t57dD+9g3QZdX6HgnI8aJblRMHrSpn41qfJ7DqvaguYeckfLN6sTcplokRA
RzVWovZaz4OIxf1qQcMp6TwYFH1Ln6k3ATQjg5/eV06xF+JdUz56QUC+xnGXf1VKrMMvN/Bv+dAT
Z1OC5AFbnAoaG1V2NyiMjyDJ8r06YoDYedp8tOYvawUyqZ19PXmBTYqSiuSnaEBL63phXiAOjxma
VhLDG1PzkXnlmia6XMhvnR+wy5Nhi5MTKt4FoOOQdKRtyWXsXzdBK06FSpcyDX6hEaG4XCd6ZSWI
4+UIuURcKpEgxXaovpLg+HGsFDq5oFx6v7k/4SZjLRclxtjbiso1OnrihfDwtcD1+bM+/PQbo8tJ
9JXIiVYMXssTtItQn5bDJaBiBPsFruoOWGMAyJjl9TbDfSIexbGOxVCorUy9nW9cJduHfPYIzPGd
a/ofo5iuIwMuTC9V8uwVUVkggVsLw+tVsCxcTaQpyiKHQuvpQGgZlSUkn7Y1LadZoy/JEvYNh0oq
iGIvhP1Eh1Sdk18wGYj9xVMa5OvRwh3DuCpmgmih8LvxLG4UOHwXlzVGA+cNy9zw7ncpyNu/+hEd
EL5UHO7wJydepatOiGig+t3gTky28n76pLbuLB34gVOQUP0TVO1AZLbfYDOqlDw17/0zAofQ8hx0
gzVm33/wjiRiA0BH2GagQecUunuT1J3T1ogGAc197EDEkBQ8Z2czndstQu2t2IfpqKiZ9PWouKhY
g4uGbeE9f3IJ2uu5uHwFTx5TzmXT75l4GlCqxbNLcjQKWuRoucn1sWjb21qnF252DQv1vxiia6C+
KTLJaUfzS7L+WyRKBlyn81RaWsfceRD7AIj8eTUR2PblB8LKat9EB2/u9DXqrO5Brh6HtsmfKr/8
cvO7VtJOZdflvKZN7AeIRQeHcD1R8V4O+riTSTaW02O4xjODXlpSQfn7e7Hyxb1NU/9jJYg00SS4
8cl7em/uqu2Qs/WRHoiC/ZWE7bpXb56C/5xSgjgf85Ue9cAUyG8IZ/y7elcZGg5vm8Vm4BtQ9VYD
hxAsHuhzAktPTlM6/5blka6SD1EMBbCX3dFW8dwDMkGP3fAZ0G3R1/WYl2t7RqPX6s0QkP2f3xND
xP/YW0hQ7fN+phZGd9SDdvwKt7shmF+cGmLMQL1XeRYxjktveqGFB1tYYiE9YhqV831A/cNQeDu3
g5mMzR+VgQmznUYFe4nPkoJ4pWq8IVb4TOGFSSrnXBlwTBpTv55bhg2C8/uXgG3TKDv9Ra5AdsDr
NyGpcUvPBvk2HDqLTic3wkmeZHifNzQRiYAnfXL0Gmvj4PBhFhf0ke7rmgWZhpXE4xavSLf/LU0F
0rK3UjllMtvx3qWeVTsHzoA9xhBWOJqCI04Q/eyx/y38ibkFai7St+N4avhyvof55JQkUhs3yqPv
Grh8OQQEfFNc+/UdHX8gIB2oEwxYgVu4NqYJBoupUTkzXy/DjRG8NKoZjQJVK7DgBE44ZFq1WqeC
F7ltuwrir1VlAuOGG6ra9WDgOgBjpZqUGmcZzf5W7ohvrsZ9aULS+TCMe3ZCBT9Gadjoqwe+RrvP
lKPpLV41wjJ6/8bPNq1VD1bRGpcwetgpoG02B9HxalFFFyasbDAmWL6wiNzTIIWhElKqwMspIHuH
w7a+P+oAihA6PyKtkH6zt1UjwELZ1VhXl1GyHShHTiNaKU7bWbJ1GapPOk3sYKyYKBIIh3MWAvW6
s8lAxhhZ73hYv2otvmun3zBuOEI/4ySCUONLDAxNbpsLH8lx24JY+Kd7TFCew5H/wQwhEu5Dvj0v
i91yB8gxwdOrLwlWt7UpPgaok4dX/0QWRSCBVeMFbXMotQJockn1KRm8+Q9wHlhf8nD18H9MNTpg
nvGsGFomOYjnw6ylmesK3squJOSmvVW5yQRDk4HfJMOGcmPSmd90Dp7Ju7DBEEXd/RSru8KXbQ2u
4wdK7LxcZ3wGHrOH2PmjUFsfeTcgbNrXdHgi4zDv7eZHjujhLdw3GcgT5HwnCoHaJ6gnwS0R4qD8
0+pnmqiR0r3QvrziWKTN+juY6SMY9RcpY5nS/lqp5coiuZeP1LGmEu7IfNahmOpDgBRJTqeH1wcg
AqeYGvnKcNKB88/YMmTPlIIktXSdEQw/rpaYSt+1XqbIEL+MoT4NLFAE19HPq3UgkKSue2sHpo3k
UMOQtn7hUi7X/mUir+ZZY7T0CUez7doiJLPJ83pO8oWTTEewgcTd824kdNxo+Wh4mNqO9snqYLzt
Zl+jGiJnu6PXu04Y+ouj/lTVXGblGA9K9aW1LMAzTbBBtJU9h1qwkjr2exU6c3g5PLc+1ugbbVMN
07tKp45Mi6y+gK/AB8gYF/AEUT/sabhX4ebICGRrrd6qFeKbm15cyjJdBVMj26k9y3ZXH7GwodaF
s4UVWInfwIMC/QDFZ6pncoqhUlXSn8Z58eSBg82xZCh9u29jLZ/+71HMBMqb27dZfikfWrLmz6X6
o85BS256YP92ONW4LXzLpLD2GQLFGoxyNm9asKjgjy0hiplhKZiHtXclRiGFIZHSOkeIj1f9FE4f
MuFzdUovlGHQV4HN9BRkRVFqdU3rj6M0ZnogNuqIq5d+Kq1wIzsiy0qAqBun/zXeW7+FqyCIg8cn
OGyoudrhHJhQlaagjSFBWsCQgTVGJ0P8/1ZHLkf4H9q5IJSRisbjRtxsP9MTx+6fvbCG+Z5/Tmg7
R5e3FiwdFrvaHFZLVIcq0EzhB0b49x6YxhWTMtZrPJkbpqT9HRPCBVrcpW+Z3gLFgVXcSn+8gkFj
HA+zdHRt1kmCXsHGi8Fert8B1cPNlZ/cvDwp5hmCV4JxrVk5f7lcu5Ka3D5dLtkTXt0Fx9RADgIZ
pvrGXEnVelTMwU71/CGziTBRNvS9bMpMAgUBTkNpFm18b01A8FrhfBTlUlNRhA8+w4VZgeIg7mEq
jUYlDY3b2+AdKtw3gYmkow2BJdxG7WElp8S1iLUy8zcA8F1CTVbba3H1YZJhkOWimxXhUngB6DhE
Z9hKyECjzTU1MnIddN/THnzR4HCHWKDf9C6MXdhhPg7fLlTdGlQPXIBq5xN8HNyXuRbLR1A+DsfX
q8eI2essQiLsYTQD9iDccYcDcJh0HLH4UtY09uTlzKtzNhbETysgASCSFjXGEngfzuUoWDZhoBq5
J0K2oBQ8XWjOd74mVIWE31bwUEjhQJaJpbnE3pqvI6fH01lj5IHj6HVGsHgMFwnvegrCnUt2r1/T
tL52wbCbBcfn0E6h8TCzLOZd3SgLwIILkt1RCIFqxdp/MgmMUF48S7ktO7nkshZVTFhfDZhC4YRE
uiIHAjuUluVWRNFMat5Q6MLQJL8TDj2M9dtQ4BKtcf2I2On1QO1qW6pOtW0R5OyD81msQKPbUsSx
tUxM5VN99CgyLVDbF8IQmeZBQf+v7Y9FqkYLTpvTVpmGPXquNWboSp9w2NjPJaPcfOuBHpT0VVWS
a6rrWR1MUIHo9Pub024Qcw4xnVRd+jUy72UvBiX//8LGTYXahG+RDlGZUKQjUjspVrJe31DtxaG1
7qagTtsuaY2P4OztKmzrOY8xbvXaTbZu8WJyPt8MBuTopdDT4FXmhz6vnJRsla+jAA8aEXqbie0h
Ak630AbJdesOarlwwBHdWdhhX81vdrTuG1Achy4dB1RshoOLTLu6kemJB24iJuXq+Q76Unf6vHAF
ncl4KweUsdYNvFFTTFO8zlKhDwt9wAEGASrwOVg7CYuK+hBGboIGZ8Iy69LBa/RyE/1xI2x2Av5c
yW44gwUmhH1OXV8Uo3VNwfcXeB6OwFMOsWUCKBmnSEzeI2j5XqRiRtk7c0mvtBEksLuUOokMBU/S
icXjG+YYt9OVETaic+nlZyQW5Em1Eku4vux2A10bTcRcAFrEDi1KjvSpz6GVWc8JzkU8hI9DroaO
EOWo2r0iE0Aibo0aSo3CGotfpaKrG/VcqmXatXeBWuLS3AM3fD69pfAwDdRm2sEK/UbN7hUQAHvX
PZzXlJQT1LxkAmXr2w+yHZClbNGaK3CwY/uIL4G1IaCt0yAS4WLWJcHF+oXtAKUXBWzbnf3/z/O+
eel8pfySdIjYyK21Fn3tnRh9ziOIz9k5JqgFY8O8I2lgPOmvsSW6g1BYg7mx3wS+aBnuYfXJgl1J
G91CKWT0R/FE0lflL40CTEs8GKiSVrjBUnTrU/6hyLf0/92fxcyUJRG/VHCJ5qrUJT8945DwlOpo
Zz5Z23JW+zhro+/GusZlZNigV2N2WqPMGkCZCS5zEpkxDPmjv7/+YB3LQYvEYsjqj8oOvmiN3mTC
9bNWQJ7oLxonAtOKrkaAOzF4WyMelIOTZpcs9RXqxnatOtHeDcuTx0xohvOKWzBvLBrGEOHaYfUx
ljUEXhT6XqTZrkmCxny+4dVdYRYDLzzUuzf+ltj2kstQ4SwgpIg4Stw/xHEe7+Q+F/eXHsIx+rsn
s+ANhkbLencWK4sAbvLFlUo7m5hipgn/IOcj8Q/NFE5lJtjNPnVXjizm8qwj1Lt7lx/E0fjvnhpP
Vq8MVHKzKzfXNIjw/gc1ESgqVDumO8WhLJVeiwK0v5yN4CicWU101De0diN3Yq2WcJtMmFvFtkF6
Mj5sFxYmIPZ7b0mVSaA0UzbAe3770IAgvuPuYwhMMBqUFQF4443J6tu9IbhDcj2e/P89H66fKtAA
txCQKXWwXcY2MsDUnxVnoVS37EaG9OD7zNcv7GxjT9bP2F3y7U1/4TTXPZ8jZXNKNqcxxeKDWj7j
7qwk4373Ik4Tt4xNriqyPQMoSny3u9jYGey5PCC+i/OgG4z+lHVwiwK74OFEvT35Qwx8vfgL5fZl
wm39habgcKHnSGWwKew2k+VGMRDBQjtfVcPrgxY+lYlON6kgE48M94WCD4DwgU+I3BlSO83lAVMz
GnfRlQefb9vblF8BYr3/q+wgDPqZQsDGm9gaa28V+dWngGJJLo2Q/QvxGLwkSYa3txpUTtBagKWF
gf+QgG03jjOI/QfbJJop18Tb3nsZIhoSO94ByPlPqGJSHBKzI9u5Rn/nNul5V20xPnROAIhEPCD4
O2rKCyG7GTRYfWJ+jmQFeeEH5acJZM0aUbe5/xlFmDcbQLYbulOKJeQfEGLMjPNWbnQqBmB+5QUD
CoTygqoZSIoTxSRSE9yd2P3ZDJEDC8O2wl8tVqCBZnLmF0QavDzuHmQPMuNMuF53DjL6loEjuGSX
TiZ/Ml9O8FwD9IE16DqjDNw6LG/c2TX3j7D9eXjONXaioe5hpfwptMoxhqm7Xm2ehHNK1NEtH8LJ
zKkwDp+e3+4PXudBzCotdx9YahYojMhkzFLrQM9GM9cIRbqyfvMTxYvZhrGqX5Ywwj2MvLkUQbLq
RZiVwhXkEwVQ9jFDuMpVD2Sfue4f1Z711YtPJOq3OfjfUZe5obi21sOz3fiF5P4rkZZvPTze7lvs
uLffQ9ZEo/iT6P8Vj/36Lepi3B+YU08hjpg3tJZWw/2NEOOa2v4Oap1LCO5bPVuefTenRkohYLCv
VH4iWy9Ba4BRhsnFzN8T8erzTxaWeND8f3YCMtoY0c4d6sWp5q7bpRWTqGYgh6dkUkZrPFW9/dij
entCq09FhccIzE+sasKhDY2mZatHFJG2FMKacK3l8njgm+7pyPD9LwEOcfKK/r5O0U1tkQhSgvBc
H7OR/aFbUHXlzj6RY38k4fJ+qt35uPCJIDNvpfag9eXdbTqDxOGmvSIsyl1b1z2FruL0Yevs6NMP
+RQcMivw4Q5GopOiuT9noQTdnsDKyoMIUYW+adxqdqhGE1qnPLS7kX9mlrW9RZQVdpU6VJJ6H7zl
+fbb1fXfvjXANly2eHjX1n7Hk/QGrhB4fnBXMDm9Ap930mTjex5LtoB8AOV3qLSrByHZF56e8j4t
oxuD1WixOTlEOVq2aY4C6TT3GwUwytXH8WovYpfIXkxo7xU+mRKMYk4eF70sHUBLsiP5bojeBjbG
cP/s7eirxPPbgtsAHQM6Eugakpae7NM+ONzA9DaLtuRl1n/nMS6jkg30jjlcYjM7terOdNkuvDkC
Rc+En+LEwI/WqvXnlgYn72ahm+IuLU3kWkkMH6VKqQVkcHSYUjviSuCMI5fQDNzrvYcFsahZyE16
AMpMqJ3ij/8mwvEAjggRNWZ7WZNJ5L3CltjvCvK/vk8pFO364ulR62LlAQqJK3pAO+1VWfp1FTj0
DZMbnBrc1H+98MASDdzzqJ2mtpdHob9vkIvrmVohJsoaCZRsuZtd9p765mrDt7gRAMH5/5vHSNR7
sL4siCXuNvKFY2iwZ9FM6hIA8LV9yC/zwp567xDiF9R2+XB+6KY8VWXu6l8YGfnA9IjKTJZYLXJh
hI7U4PtdBXYC18sNthMWfOmfLZkoWlrwmpmw5uEJ8Y+i7A6+Q65E9fjuFgTg5+deycJasjmcL0Gc
ngN7QbvJ/bxRZnShlINLNtE3Qbg5eKRt4ziKmtus4Z/Pw7lHsm2wWn6NKLJzSYVKq3NmlcXee4Om
w83bmGYLgdYEJr7t3HVlIdqar4xKc4Cz0Ts8ihC0T3xushf/0ByJBosaMZ1GTJhMCTUVvofBIGkj
gjkthneYatn11Dh5owgwO6voQAF9jsz/vVWOy9dKuYCYZamox2d08m9oNxcs9Ay4aZQ+RWEmeqIL
+PEHCjMh5uriRK5yIZIP52LuEQskcJ49pHmydAU/T1S+M3hpJPVnTGejrr3fMWkrbdiP05NhHmS3
sxyf35dxY8Dbktxq9mnXMKbOiF8+XR3BRwMM+Xeij+dI7UrjiQYEkeJtna5oJz/xMdkxjiXPiT+f
wj7LhK4nsaAKtjWcWuC2ihaB4N4AvxhMrfTSoDlawNto5m14t54CCXSuqexjvHY0v7ytQfyBNHBW
3KoSvovNY4hQ6H9y/4s7RT7dseIZ2S5JJhrzQG0b3BtxsYF/lTA7g86oNMHlnXtRAV5weFlLXQw+
lAMnnRC43aosV9H1SlYWZ29Z92P1Sr92GMT1lNfwEzV6skaZX3se35Qz8IIZv504jXXDd8f/xlwf
Wm/g7nBa8eD2goi3uEBQKte/CfcXu/a/vWWhQb2Y0OuNCvygx5NYnGujRI/WRjUfmdOU6nqD5+0M
AMoCQvq7Jo0fVUSg+uA4VI1sesFl3I49DGalMc0dUnMOdTT4b8GCCakYYYzz5WKuUsAo/0+lTJ5e
VHdDEoX3aDioCGffkrWe6cp8hrseLw8/+9hH53wAMZ46KISfpYALp+xItqnSUFc0C1H7gv1TJten
goqwfXFCRNm3qNBo95EtUZiagJvSDaVr5y24Sapdfi1Leg0hCpcwuR3yocfpoyw3/XHh19QFKw2w
M8saVgzcEqmav77ufMtc0fL9/S3o9qEt3SQLHwBK8s/zzE2XC4oDXnjFlw8v9VhmIkLddO/RTu0w
jyA5T7MqyktMLkiVZAUkoEOVnOyTzZVyuA4ZDW+ogRB6sx5CLBtDbsv5/cBG7ZApBX1ILAdxpi+0
JUQYo68vDxPQbjmNwFTcRO12NBVrABv8Tdn2rgEyUO1WVrV8Afrxq6T5MIzlt8ed8qUgIatoAV6e
b3q+lDPiqYwkxg6Om40DY5DxKZ7oo0uPRSdGeKnbEIpfVrrVEcA113QBco4sZ+sGs9rI8CaRUXpj
6Uy2mNnVYSoEV2Ju1wbz1IbunToBh3yQ5T+Pgrvp7mrTEC7BeGFLLR6Ubpg6DIv2dDGExVpJHgNa
L2G9UIeRHyG/trc4CU5f/EeFQAXOB8W8zv5ks9q7Oj05emV6Vv5EBFAqkIZE5eDD8Lqsn9PRVp9i
OMACky5lEiMLvSYxZi4/JscooEisoJfe9U9ArSEK0Vmi7YZzbkAND/M7ePKJ7SDe8tqF3b3ExIOQ
waH40hBjXUbx33vEur84L6Z1L8PajISa/2pBldSKXjJRZm6va4lESW0B0e8xGKEoKkdlUgBPJbqu
E0763rfzQA20oz8DQ5SROp88dxuc8zI3P7qFamcouo2DYY/Pod2u3QbkbhEphLXs7psJUg6Yz/tC
4LomlVLXpAhg7VEY1TJQ3r/ZhUZTnOD//p7M2biqlyWxBCo7AUF64yFgr3siEu0T6leLlp1NaGbe
SM/wm22uf+vqyOsaYROyTFCSXxvsV+YA8ruV0ddCYubj55T7xbHUmNBGpOvLgBaosUmxroCBIALP
GrC/8ovl+rhvdsC8Ro4lR+HIWIsBXlTNjar3+0t/TbDOeW5m27Ik+Aa37IETdYIeVyrnGjZ+z8GZ
BrovCv3f6JkMdLlN/3X/iaRWBcutyupJSEZ1rDHw2EAo9Gj3LXMI//eVtaaV9bABv0VxPSonbJLH
CA5Cqd/nrCCqPL0nmdrL5d1DUwfSCzwdIbt7C0xjoZRJk9OC/1ysC0AKmQNkCGg4NXuc/usaoAR+
12+yYy9xkzPHo3WGEAEpnXs1XNFoE7Ey0iolQo+nLdUvjlYV4ofv53fcwBkwVqtzR6fVedZ3Ogb4
WBHK3NH4QuoW4UNaLqt2J5yR5g4TMMO9EMXBDpiAgvoX8NOgkx1tFUjMg2tLvcW+Fgd1hGwxS5bs
bFceoNsJbjy+D4pd5+J83yibSzrkjzqUw2tx8fevA+mFK2Q2KnDG57oL33PWfpyr3396HxJEcjIf
CmlTV09N0jRkOURX8iX70qC4CqM4QFJrkC0dWuiu9SNBxM0QVjYj8mYlwfNNRj+hX1aMT5xd0SFA
of7gFNKx+RrM0SbKfl3rAR0MhMTCycsj8239YUDzAOHs82/6MSz7tiY+w7j/JDQ2CLHNIaiTXUWt
7kzVw3cTF+mpsI6/b2WGaFXlMP6FzH5ys4ACCBtoHCtvASxqkbmoHRXQhjIX22FYmd5vEFIXhySv
1MgQd49OEIuOOGEzaNTF7g6XvkideXqFjZY9HnJEKx2ZBeSV7wYlj4UfHkdNJwJo0qZrPAW93eM3
AoO+H3kwsL8tL836EG2wL87TyLtgflktvyActzYcjF8uTitNNmh+ZL2b8gtCTyTTeM/zK8tLKe/P
91Zy3ZJVw02nLU1PhnZIDF0qP/m7EjLV0MeM/mXHtXtq7SRZAIv1aC1RXVO2iI/RbdNKs5kjmbeV
IrQ50mbEGg5/tESfps8J/hKjuDuq1C1agoE2mgYyDymiU1MQYAsyoVFDtKzmp2KC42SvwfXoeGTr
Ydai2SruobkP5yZ9Gb8eL157MUm1Cp9ezWpn0DqGJ6olK/WVwyMolxrhYFEkQjDmZ3FWODZrmZnT
qo6HGubCtfQcQ5CJofZYoLYSbbs57l5mxcA/XCzR+t3f/PqoeaCeCmT7LI7QSr5fPSHCXQXYMFD8
F59piOw8p6SCaHAsM9id17S7mBY/HPv+/h5A182ZPbqaI712XvOCiLqSrSicz/M6awebAnubjPUu
JGAiNqBDcNzayVdKze2BoYtL/xTsWaMbgTcHvUJ3Rj+vHrV4+hCXeEOEdlCN9dlGh2lXTUJM8JIy
4woN8lqk8tykHFUSfeAE70lWFUzym69g2xUXXbx4YgZiqEgULnRpHq3QM7WsdN2NX+Ud533v76ZA
wlzugw2tpv0nOrK8GDQeiPbuqogRyDdLuFhITVez2Xx/oc1npzHrf5enddLj0hleWa/Iix+GFiJE
uy1AfpaxOofRZE4PAr4xBy5RQG3sswKsFPX1cM6HaFEb7puTdU4JzN8++hJu6cS42RQFnNGo+MKK
GXOIOEuaXDPE/Qh/Lz8BaMNPvkuZfRGZ9MrlPFZR3YtmTjlOtjD4wIOuCiM22OcOta4h/I/YFwIh
FyHzpLHV1FGXh9eZZDt8/2pVKKdb+b/s3Ezc3vmJjv8PW3y8HDhbxlEDYVOHpABCvr7/V3HPxgJ5
4zWFaoSYmQxj/7izC8PmrLvh1PanN9Bi+zNMlz60ghgU5za+JsftYAx446yDtBTteRuw6l8OIlk6
dKBUZUGeTvOrJWuzxh1DcR0Q6swcpZgsa0VqSpoKQ5ImcGVv6VRabsLyZdw+gZm3Umsl0euN+pnR
eN6v0ZhHIv3PyRZn60JFkmwI4bGwGvI3PbSv3QFTQRColQdNvn4FAEXy6qIZnRHQ/j6BEWQbVun8
p+F0dPS1d26AJoUJ1CTGrvG04cz8upVKnx8SNppfvrD13AO7E71S9qIb0Z0CFp9nDD6eJSgy5qSW
YvSQeJycgjqHAkNYahFksIE6+wf1YJ7JWu4lh4iSW1hTb8Y+E3rlIMfGghEdp2ZWZN8+yB+phWqz
I7fYzmWuKhi5RPDV2KgP0wmCfb3movn28rnfEW+hPUPwxdy5LuFcqUNPcj1umCwqaYDwYR/kyOCp
HPGfRXyK49riEC+D1l+kszj7xk5cSN09An3wl1qM39UZEbsTN5EyNEoWurbdigkPJHFIn3l90h5v
pvvpWdV74vpQd1IftGn8wc4k40M3fo0UsrxzsjfQqDt/Y0iz0oOfrxCqO+5UhI2vhu0Nw4MOX0sM
/WtBPy6un7cbiZvqsMXGwZ8Xmz4k6nBkUe/eA3p4SgVupqT1RAJWSWqA10uiELZO+VDdkVTCEUHR
2WkOJmdwMEUf32HliRBc2tvvhWGGnWC43lkYgJr5rsxiloEilIZQf/gfnOEOLVaKJbf/gToxoT88
jJLLixaODQTiWefgboEPcP+WQJk+95Sk27OeNeGiL1Fi+IgMTHTg6GfKvo4vhSdlcWudOnImOItT
izmcVs3iGlgTsCxLHFDwc4djWDOeBQdy59S4utCiod6uJwdJngb710iNmr4raUf9mFe/G96jNRIa
hnA/UVGdnx8MUnDKOyYeREsBWcoaXv2Y1nVMG6sEwmU/O0fIomkse2XKoWkzdLHB9xOKqqoSi3pI
+HqbnYYSNvmk45ZRDaHD1zSxfGDN8BOl04MAnCWbLoT/I2mHMydxDDZu20DcM36oHd9MpxZueGud
q96X5ArqgGv5JeIezbVUppsTTUTy9wfB+DWQrxkOnEttdDideZiXuZGp4Poggz1LbUBfgTQ9EZSH
3E0d7MxOMHmH4jJxM5matPfHheEwQP6IRvTQMoTPobvZSaNYuUbjYFvBgQi500I4naegwTqumj2E
SYsp1h+IqM3UvtuMEo4jDQAB85pfEBsmRPrRKXBUTWNNw+YyxCKE3+Y8tm9z0jPzYlF0ikT0LUON
pcXWhtRzJf46sr7FzRvfvCS1jp5mZubsU3plbxqnYVDmYz76F2Q8//4viW2/5ROrWFzeok0y29P6
6xlNYZ0IX/nPPKQjeh1sU9IeaAfC2BA9B1rdoy51P1qJSJGX3WKNHwvq8HEapNrHZV2KTuo3jwf9
kpHEurhu3lJLl4HNy/nn9FfIA+1fSJkWbbDjixE9y/w4O9NDVIAY6FMjID4sMtHPeF38KZ0eZDRf
BWHKVRHkXy1ip+121CJehdfSw12XaVN/kCHlXI6+oLIoNit2XFPcG5lxJjMCq4W5nhaEiwfSTSYL
FOARm/jTalCQNbRJj3XbyklXbGWaT/wLWXHkcYuvd3BTDZsXv88cIannWaMhbBBgG1QxRr/rO0Z/
PulAF+C5Cipw2M4gjcOL88GceZNgmgOkiU59DDo5af4Ux0GMrJEwPcMUxEF3WH86ZlPfpubl4OQ6
Q6eo/io4NHQoUaMRqPrqjaa4M3hA8iihKWHrAoP7kK8PxPYRtkaAhcLV2g+OraDrHSeTglE+FUAr
UjC0umnq/sY6Yx/Yqi+xKuJNgs1TDL2ovRhrwLg1RifhNG1bk9L1RNcCqLwykZq4TfqZsZOMJhvl
DoMxyU2RK4K2oKrT4XieDBM9aDhGx5S/jW7F5kcvSD7mQqmVPpRM8gSQDScMrEob4NeDInc4u0JQ
WMpm7LGhTIKA+GCfQmimRKwocJNq8H7wen1yVUpevBMh+s+/sMmpG+f4N1zvti3omAEtI/ns45Sg
MUGyxXEetY3Fo9vP7XQiZ3N7RfdAwclLIqx+cdmO6z6+PTAyrVX9PSQXU8xtul01CV6CU9MuNTAS
FZtDgU5bwRfMkya27VewlJS1nhbGDxnSIFBYbxCMs8RzsducId3X4tk40sm/ptg+1q2SfdwMWRY+
HpTtk5jiadr5hEVZipyJ5rgdLL3aJ/o0zbD1MiZMka/kNu9pxkBGgL/TPIkYnuZ9Jd3UakOio+b3
5X1wiJCrmCLJW7/ILOtT0Sj00Is41xAwyTA6hLwy+akwcwRbXKzuLXacyKD6aLF8lCAlY6UGMa9l
4ya0SZ+yLFZrCwYI+2bekCoy6slxS7EzR9oOqitvMBaLDfEv+HyjURyTawEtlCYfOuZ0UIJSBikd
ffc4jEWiTn/nnfEJy1F+eqAyrnCdipOjEYHNQeW0lD8z6G9iMO7PB8LNqyXn4ef6O73PTpr57Omc
7LsDlODOaR3wkHYmUM9OTY+7b6W0PdOQrJ6YLwvth9nfiXEeZ0ikHzwpsFe9OqrmjgU2ORg4zX2b
b8FMKQ6cTNM5idD9clms5XDgZPX+kRH0iaHqBP02awl+bgFjYYqZ4McAWQwea+P+L+9lmf2Ui77n
X/EOo54Waktv2y2ieW81EY6uVnPfjHRXTM5GtO9fnRDx5nrtPXvrDLVFq79zUpy1MfIF1TvpJt0N
SK76gXiT8BKoh6WoKkGF78mLTS4ltDVDeuJLqSd8sGXdmrDAiGPwuybwg5xy/XVaqtQHD5Qt3ajp
xyeniMF/lu1vQrcG9asyMWzHgy94y7Jd5s9QdrGWHOJHIZPYOy9Pi/iKdOMJT7ZudfcGw18fKnZZ
yMlOdCg9eOlZA0jWfpW1tubUk5gAKEGMuxFhkT25hdDk855gnujvDLdENi/Y1XKONXDS59s/sc8P
jJv6TCddrLcmOsSJmWGKy9OpnO2e67tSVFNBv6OLs18B7cqy9iLmxYQ2Wa0gM6kORo2f/Z3MM1et
oGkCwTc3TvAYmoE6LNF1z+qccVpgmNx8X+G/tkuKjhTRbfMQlVVfpDZt7uql/8H5pcp51akG50AS
nm5F+poImSPNtXMHop95P74Q9hJKGr8iUY5rJkfL0M/BWkhOtHn48M+5Sm5IyzkPXmF+zUDCvSF3
hBVZma55UUk2fxCbv1T+2ekrIUkA3urXqQjKYhmhALUFXR8hIg2LHudg7Fmz24jpH+s4zbeR8xHU
KcsjvkSiZz5vAtREP3O94iHT+p9Ow/qQIO0Cth+hnnmR2YO2RW5Nyel2sRsuw9YRdCLpP08f34mV
sgnOnTiEDTbSDLG2eoNyflC2TP2TjSGWLRd6/3LscS8Fr3Mvr/BqfnKvEXzWcK3GKcQ9NSzFtC8A
QGQFPFXODHx0+dYmLBJ9itf7dmj62w1eju1KOoelyj0V99+7S1Wo1yO50I8Z6VHbQCn9XoKOml0O
1JF+YFUJ3Z+5cyHefBLCOWEFZg9ISkTKnVEUAwWC3dUpQENGv7qjTg0PgeGLELQnGszXqLNZD3jm
fbCxbxghdj00x/YbpOTXAXc+STkWL1eU5Wl5teqsv6Miqw/QlAtniZgn61VCn/3M55Vg8I/At7Rb
1KSvkReE+pnyNN2jX/qmBowdHTKINWjwbSfA956fWbWeklUKIpOJjUhftTaQcMGqWiykrlTb5QSY
TKhgWVT2wQXIDUlqRgDrBlm1t+AA5kifEaHPjrMuWxkuFO0LBfK29ga5lisFJGnoMOapFqDztOqc
kbha9PWg5EiR3Yp9Sk8TEJYaR1tv4RDq1yhtLgL4x8xB09u4d7VSKu8EMULFM8lBelIFz3UNHj/D
apU1sZO/lAHSUWRhyNCWrgj/nOA4FsOcg5XY1XSarqGWI8KwNWE0UeYYyuuW47+OKpNFddHZJ6jF
rUuxu1EhZghDG/kzoGVMIrdhxXXsqK05HixlofYYYYiF+PQZzH8cmhOPkkgl7S6mNhZakKp8D9Ks
7dbEZ8Q/J/2kPCXAaAjnRg/hUgo1iOs9w4x++/VhzC38K9bJ0/u0WGsWdhUF9V5IKLZe8aAmsaLO
NV3k4BJ7a6z/xVX89tzMva1AGbH3MEaeWQrWSx2VBscY9e9HknI2QBYQK+30LokkYdvfucqxUV2L
BLme4vyQqDn9Pqm5GOdoqW1Bh+PIZpciRjd7BdLe+JmNsDr9kVh3mCK1nqOjJ/AaV8zRmFYlCKWE
NDSU4D1NTPf9//Ls3YKsZhNr/7UavGcD8cIr44tJqO8Z9CUm2IY881ke1AXphlpq6LuZ1Df6ZEEN
/0Z/3cJPaoNqh6gbVeMas4UKB0QPolKnXBAZEc3SZg9YuhulQuH6oN7XZGWUBxr4TgLw5k7lW9tk
QVibIm+QhtqbrWq/RzK4uCGAh3vmA2tm5SA0h2de/m6GxIc99t/fA9W/2to04dPoYogyMCPhSJ9f
5a+FBGD53ibmTslFQot2fMWrS4mcbxf8Eui3FZ+umyUDiSIS80gHYAIQ5qToqNP7EJlXPDhx59vI
dtZ7EgkAhS/1vQcbRrxgTtoLH11MRNeAIQulTUznH5NMh5XGm4J5ucYzrM3QgtTTpEpL5GCIfAMn
Jfyi9qKN7vnZKkmHybjaJL3VgqiIBP5uxad0xuYcIRN13A+yciUeyCG/NfdsciL9SabxOp8iaWSm
7HF6c3uc9e7DssdTOfpcLRr6zemQS5B0ACgqLkkwn4J0SBRT2OrgDouFrljrhin37PTX7An3Xq0P
cUhFBhDf1Gc38Enn1P75FAi/SGMsJ3YpLIXjaqD3b0fZhjjTZn5IXosJArmTXhKfR+q3jF81dRN+
KLQhdFzlkiELf1BrTyxZeRCgEg21Cg0BZIp7EK1xcErdyIK9Z62nlG1elKn9lb2xiECuj9TUEk29
Lk2H+YQCwBvhyIIeJ5Y+gQ7+NLlZ7QEknrTM7RnqRlSmcZs1dG6VPO7pLD+9K28SiE2fJ9VmSo6O
+fgBnLqPaH6PKADqjQQsC0l5c9nwyffJfDyfCySwjEXWgAjygmZui06WaP/RYp4WzifyOTn11K4q
94iYfSvRu3PtZT/H+Pxz3mP6o3gkO44OZSqVWgmIr/Bzw8S+M7qbXeDsoJWvqfGQiwUtuhAJWIVk
wkJ8ArVM6ZuTDSFgFDx6focuNx4gR56o0hx7cd6YQ9BWmq9DymeoIpL1ReLNKLp8IdfYCuimfrIn
jLt01O77AB9f5/Y7J0ttMrPcuS3bAdNgtygs1c/wu+ALIi7X3zKEr2LbmWuYD/kBkLwyAVk8mETT
MI9XZdGyGVpIvl9kMGphKQZBpEHtWycEQRSfwMzKhxootZ9FJy3Tyw8DeCMq54dFy/JGgvpXsQ9r
YqsnBuYw3VfmCaCS8QYeN2giH62GwJoH6SupI7sT4gNk50WS0Q2zQsP57sbaKrtdDLNTj3TADSHl
JMGjm8fHkcpd7eFXh9GVI9ueBj7dUq44MotPeHfwd47c9pTeq6jFYIP4zB1gKNde29lOWCDae70e
eeS1rV/YSrwpQvIvE2LD45Aw3vqbaOF76la3ei3nlUDSKfTotphkJmqOzOFgH2z3l8yGNivT39/b
yPImzXOfjS3zEfFqldmogzNy7oz9snIT2mc2HJ14sdWW4U7X90LVo1N9gvXXdNb2ymWHbXUWIUxX
8J4d3HIqlA99Nfz/OdWq8JTIuB2izXbYRDn5lYeLTn1OJo02VePaKFjO1m2CGUXCUnNpF18hWAcN
FtDGZtcTdTptb6uu3BKn4vB0GA0cRoqUQdrIowN4b2r578ZzCPf6qB8qb0Wyu3Q+vgAozBbooAHt
CPLsrWHubbz2+GoYn+chuYhoHU/JXMx6m5XqEY/Lx+p7v9nF7S7etgkm3ZFgVbH89gfIs3ImlC6C
1aOTFN9Ad5XbwPLMozWkiTcbOr+XO8JIMer2HrKud/inbP4CxvKAkR8zQIkTNAv7aPWmwoEVtq2O
MPxKBDPCrlJSb0WvtpfAsNewI9uP0MzICaJfkxI83DB5HDgK40Bax3XitAzhmORAMR3AB6+cj7SC
5I3wZKfGVkg3YlI/hvM75iaKDEfJN8NlUUPm2O8YdJ8SPaKcp8vYLi43YJMhTZcIgEKnrUOx6fWj
n5wOhC/KnGZuLz0CtDPHAxy+iQ/EaNJN7JkQA/31x88jE0GGF6N1zT0TW4xNVMQCGlAz3C4bjN2z
zOY5QjHy3bdoaWNaOf/ApzG7oTSA7QLIHTcVEwfNpJFDOLPzcDUtIgdZfmxppcEtvcgedVttenx9
P1J2SD7LHr9ybFBPMZvHg+Sshpa6U8QbfrtlYzljxALJDTraqJVBNDVX1qmHZvsa1vwcYk5Afi7S
dtbxBQoIoFdTjDpb72uJZueWmKY6wKtfcQqlhbjw4NHFsAtTTYUQJeZgUmKi3rzK9Sv2YY1slS6s
srsbc3AwkuaavuL1cWWYnGrzlPRdCiM4QOaXfEC8J4n8HkQGMBF0hsvT1gy+o34B9ZyZB936xAV5
cExR31zTSXYs5RyNKwK5irxlKejvnn8w1hRpAimxFKY9VB0mrL/wbCq68+RIvIM56HW/YNltnGpd
hAZ1JM37/4yFheSPZa664TxQRhF+ku0vF7OmTL5LJXtYn+/aoF8szv67RIaQK2N7KT9snwB50iAo
g8JueGSmwhJjWFyNfgd3wLqcK1NnTEiBR1FJQFdxZ9SLeK053+Mn8INbALmLgtUDVOCV385aHh/e
OPVoq2yHsQd3JjrlOOLJytNZyuxXg0PZu74+LE6ESzbRmgxS1VF8Gdww/xr6AtfIEqwlfjBVdjex
PNSnwAMcd0Dc79lBN+3bQVqOeToBDVKMbWWJXW8aT+Z7gddVhZE44KhcK9Te94VixumF95Z5FyNk
1850DeE4y8sctXTpA8fw3yZ47qQaCSdCA6Qzu10jHtwHKcXjGoGG+Jh5GsN8yZfhmTAsmuChMmvE
MDqqNExy6KXTNAnUT++rJQWSPPe/gQU99uardy47buEV4BevsB0AxG6L8gYcwA1mx+OAPqkBV89B
w7Dw81pwNK2CBmas1HE3p8Cw/m7qJDF/iftqlJFqgatQ7TNY4g9nezpt1lEu0P84citWrirywLFv
IH82TdwZOYPxL2JhTTNyjTCazPPafbxVx2nsftXCDx3vUeC8VHIZ6Ep3FMhB5ZE7+ejEN9SKM/Gj
u+95pjPZFIhfqtXdBadr7TEiIZvyKqLeCyE/ELmxrMdETeqTXp+RUc1NnUiK310FVV4BKZAJVjVs
rVQ3zhfArG5LFLnixTDSmcfHpWuGB+F7r4TLt2o455qjYGIH9NANcsw0ExKOlSmCixdJU2X8VKrf
mXRp975XJPeAlnVc13IiUVE6ECnWdDdF3O/VNOzrePwOSwhnviuaIeR+/tkfoNx6/KhejttsXTJx
b3tTbwkLSTosA6yKOu06y9QiedOydyi5KA2a7RF5iekncqKHQQqi5Fyr/U60OXfOuWBxtX45fPic
1ay/pBHtUGAWRB0of0m11m5prxxe+dMpTmwV/ap+cgw2HWt4DnfAs6HQKqe9QsatNDVpY0rGjr4g
hCHEFtl1enkF1xLdYRkUorg6gFqr4fvEYGBt+EcWi3dvpsYb7qpgA3nQXN9svQGAFuripAf075IK
Nb9suj3cjQ1sL3QMSEWX6sM6Ey28rH8N5eHWZBaZWq7HqdotBczwXfsZkSOHemQtCewdM9eWyQ7D
YiSj6CvYKMAhLaJJwCnRJnWOssASLAp6FjDXSOV/AFe11Ebw/ma5Rin7LJi3NpuDnuL1wcX130aA
OBJvhlsifHdFmlHqGmvGWAScqOYOJUCHBdRluiqOqBYKAm8RLhQALKUCItVS962jf2/n2aVpfTeO
a2P0BxdV61NhORwrGUzE3YlvO+zDqKLrcV0ge+qDLmXrGvUHp7Q5eJe7cuzRh7xEXCN6sysKQNuq
CnYTMlkVABTIcpO6AHzNLiUv78BtU+OybSCs0X4APMNU9rBhHoUJ6RbWH7EvbdI0GrPfNGS4GZv5
/p4zjrZ3jYP07DdvEl5jso9rV9pTDBzkh6p3oBPVBC2Lxj2a+U1Wbql9I++r0564PadXxbsjv0Ev
+CYrVbao4K4KBBb8i+u++m+J6ezwkDKKZyfbwu0C0qcw/zVyOz+rjY0fIblkqWvTumC5aUveAUmp
lp1r5Q5LkITHXpTNNTAiHohyn6twqtznS00V5E69FmVyJzfCOmtOHN+nP1WMdcGJRYvBMtEAgDLm
M7hfrWv3vcOBpDbEsmGUIRJgwU/CyqMBy1uu/G20FF9qdbpgYBZ9FgWC1jNQbXwVz8Pq4+rWqgtJ
9/GOxHru8JwowCVy0XNGmn8QY+7QmwM9GZQlBIdQM/OpNW5FPJcE1PKLOESDh+5pw70as/m4y5wm
zpjwAkKBGK5UUSZQgyY3cpYs1Hx3hzvVxKWIxVRuWxUwk+q/FyCrWI4aBE9i4dtNcIoeLk2taaRa
bhOHSWFLs1ndUWriZXq6jUZfdJOQJCCfKmnWq/47ZL2fugEP/93aInNc27w3gR33mRz3BDbCHbOa
t3iGPCSTa5aOz5I0eHtSAcPBuxdxoZLpeBQk8+tJuv0YY6JspXBpU6f91wBogKuD2pSxHu6EdpiD
hh0tfmNF85ZcmkHMuDQzSBzARcamggziFftIv3o8SUU5pGVOA2gOrOtX9srvbNAoyOCSsoDos11w
d0nPNyxwM5UKSDe83vgkqtQDAqi3rHUSGw4IveAe0zvKUqktOslDKIEX9UJ10xeixx347oofqJkm
xjqmCvdifxBg75eKtVHkrXfnwmsinWZwco8sOMeNQUhX9DyNfx3eppdI/n4WbtBOCNNPPhSVM9OF
F4XAazan7M3SvqzlMXNhCn4wEvzFcmM0onAvwmIuKx6caEY2CM7JoB9KhaLSk24u5y5ONhLBoqxV
tbO4mst2tuVKOz0PIGiwexZqFU0e/4u41KDSVk3mQh4sxmvpUkxvgbu+xAW+esx274sjJb4IXmCW
pCArjH3zCSHBQc5eTRYI+xNhzK9pRZgxCZM/JD/dXztiWvYUOuMKkZ9OVdbh71/JaBshswVzmcZQ
JUKx5ko9T8xvinGH2BMysLY9rfTNWF+vCwt4GhQ2B8oEjv/ovk5KYmdho0mWo/anlzWJ0juQsPcF
t0Ls88S9qsukWpHP3jUaNm0KkAsnRAd8FA3zaVkCU6JK22lrQJrx8QpkK5XYgQdYnHOAXL7FUxdp
EP+kRlLDPvMGVlxURugApT9WOhJeGWdVv/IcYO7rUl1+P3YbYtwZ3vtVDbVC3/5L3Ek+1KxwpMoh
h2wVSxoKaydMRj1cLm4ToZMDKj7Nrx30MpCfp1+2oBQleE/VGW1jXIPMlmCj/BgyApev4Gace75H
B6aZIuyFEPboTD0Y8psGbdmcJFMrXPOa4oIm0EkjOl9Cm/UsaQUec5waZwKkyETd6K81wdxad8s2
Y5ykBb0cSThlse48cf1ZCWxq3UAdDA7GvXs2ZtuNwhC4FvQLKudRYGza7M4d07Vk21Fd2iZ4pGeQ
teE2KOpG9+Dqz4vmJKLJfIgcoJQg5BqEYCB7KgL3P8cuSzu4bkIBDIs4uc6o62z+qzT2wafXlZt/
u6HUZCv6Lj8siI3U3o7THBfieayqYDWsKIOTSwSkVWC2XbrEBGT4PJqj0sc5U6pJO5ce+nY3Q/XM
qbS+jQMHlkGtk/mzR2pGPuZeJ4kXlMtAGY2L00TO7wUXrENcu34jGUav++tKluod7ywypqJo5pbV
LpD31c7SWw+bO5mtOehSfXdQhRFfSrgwEq6CedP1GbBVDQgG9l7CK/bGFYbj6IwMfbMHwjTPCuUa
zs//mj2iQ/GKe08b+AwHvwOPPY1pSV7r/DurJM0LyTorCOGiHoR5c0y/tbS/5204DOGa+QGAxl38
H70RXvEnn0Qecj7uBa7BQUy9sTNsYt3jQiOXDp9uzv1raePlK+oPyGIU3tojXtE0GZKzuTlkkpSp
eF7ufyJN9BRoNdC7iwBNucXHFOaCOC3N2QNnQK+rgUXsuEyPY/9Nv2I9Or1TwfwOQB6KFltpTNJ6
fJ0LLhkaiUxQqNJQuYrWXcNjRYEYhEvM1m+oqjPXOuWjkShgiyXkxNgCJvVSsKn15Z48XsXZ78H1
lhhzr2PtlTFAR1ChfBbJmsx52Y99xR5LzQQGNDyH8tcaZ1XjZZIgN1xND84DEhCZOM8jrFVR3QY0
nOxr13KM0/ng7ZY/NfDNEtQmWCAlM5GUDC017rbIqcU1P7MJCtlAcyNM6Lq8tDy+xq7TojAXazjR
Jwequ3skI8noAbiuB8hf8pHYyTk/Y/1sHmc1KZdqr9tDdF/N6g2koPSzNShfolb9AMSopG0ZY3YE
qxhE+nIXrshAiSosbv8OQbjqib6ULOutASzhFrt/+Ggox63tDRHu+5K8WTpl2s4uQxdEKjtdRkhr
4PO+U6bqNpiHrX1KXOniLvkGqV3hF1bXzS9Qn1aTWLFca5CpSZSyURoUG+2GqJQYoniC6DiMn2LL
mt8x/2qEHv/4Oxf73t3L9Evdao5Z+jyf/vUdy6KX41WXM99bzBzVdQEx6W0biyKIodK939ioLPho
NfMN7ouZ9hgFXZSinn3lWpiI/qUpr79mnDYW1niJ/kC4RLmNZXqu/SJqQGG+8EfOgoEBCQ0kSV3/
Lort4R+mt/Urt0uAAngGoCLmw1DlYlU/RKUXiXlYtrWeOyDyA6PNjII65aL2D0WmFHUEJNrbx5dV
2qHdEUeEItIk/OGR9NvMgS02x3QCuGEImCCtuWq8XqoMY31FQq86MHgNcPsbIFlEouLsLz7UZ3Jx
/UP23ZV1mWvITHXqSyLyDJNlf4/LZWIwRr8ZrVBcZdM8G9mZT6JOwvZsBNDc+DxCplvErtKZ1NBh
1n2wSfNk4Rsc5Bym9Rbe9+A/WxX9DqqYUDkBAdHFiY7ZSqgRaQZYEH00mgYWOOBRcDE64HUQ9hDM
FfH5Ri/JFJ5JbSvKyO6zktpgG54xHUySslJaHASt/LUA6SBiHhydEvJibqqnaDdxr/aWBkWqXLCf
m4LvOiF6nC4+ORLdTqgl+oKv7ESSYBflPaA1I+iRFjLfWw4kTtdX0Ka5X0haSShcPMSZliz+WXW6
fbQpX6yv8xUjn4732seu1u6X8jgVpHcw7xBdZctgaMXCASLZlx1Fqadsl78uppy7SRehsUNTf301
wpHKNM/wgGkzD7FrLN+b0qiKjRsC+1OLKJWU3sSg1HXl3dkhEPbft4LcrJPapGjNw/lYW5TeA7ts
wYAu0jRKP8P/M7mWUIw73yTqnDgyE6WDSCffQoZQM5SArSdvutdSevLzbvE6CVGaw2RkmNGAlO3R
rWPBETWsyA+7JX8B/nTY+GR8YY83OQNe34rT+IHNaX8tCLGbTpiIFisQuvxeJGsYg2jmcsHzs2Xv
16r9qCx+njbKbVTf/CagxqFt0+VaOzDLDyC8IJ8JaaiFtaywqPI9TYD1jgavp1ZUne6ItPEp+toP
YB5hnm82gmNHs7Vv7ZyTo4fv1m889xjY7ppOvfP0QYa6AZ0tlqaQELgoMti5iX5g5h3jvXLhNy4b
9DfnymtQc8V3kaP1swvUe3QJMWsI5v0q/8sCxw1A13MXQ6MiwrpWDX5owiO5x6/yiptE4mM6akWV
Ee+cdUrlBqD5O4fgve9b0oTdsaw4mu8YNSaz/3lLXNFSGTF3FF/Cxfgh8UPhxPnzej4QfJ4vG5gz
QowuYcn18BzL7Dc0y2GIOkated7+937f3VMOt6veyG028VmBV7Me9yIWXi+BurstWyTD6WQmQGXg
g5OV+a8AvYjHtDJpLO+b22E9edAj9GIW/3J9U7Fd7UNuTOpVeD8YCUEN/b484tbTxcxQpDQUxtDB
fXMGt+87YqJijUchL6mdyEkPi4eAOSBGosatCuGTTksu9bK9eHdaFSfcHRzYLJMOwSND1ZkbArv7
N4AY/YNYL42A7J+qdJe7T6NI5eL9SVumRlR2y71uylDtM5lHRfzY9BILbjuq0xcazy8ETUG0a/f+
iHU53D1YVOtmwY9y1m/n27mExa2ObPb0jCvIfooOzW2WDoYlpqLALvtlul45faVrmO7ZnBeYhBNe
O4lt9XaG4fBhHKWHkxuIx1bQBXzRJbE8CsxC9Zh7E4+R0raLN9Z9kPWzKPnCBmxouR7joJEuYf/N
Wz6jZAJJ14VAO8AyDKRmuRsMe910MLaMETWnSszY4VIAUugJoeCCzhz79dbh0Px8QeXAf65bfmf5
cjAYf+JkKsy6new0EhBIFcDk9FIMbhNrNf8qPMNDOvpMS6PUG881lC4iAnmtHhWacZ/dCpOcHKOv
C1FpGcXjM9zUVQ9BRsQrUtqACzU5RwksNLvzQCBwTTdwzq9hnxFDxAaOtFdODrFH6cdKiUd9lvXV
dNLI5iO0Fy/QuRWsBI2Dw/rgilGS6vP2AxLSDlbXD9sqFu7StjtLaorDNIszXwcCLL9a0nmZCyBR
v5vKe86Zmt5PttoKjYiKjgt96bLum7SL0+9lzU/AooVe6M7fzO6wJPbfUqFiG6VoRj7cdRkNy+qn
OBv/rFU3Ld1ciJd2+OZlwL49s3QFqLjAjBEfZvhYI4eHHMWRWV82GcMzZ+KZZcygs40WAPJsmmLj
iZLEQehP5d61xTWietYdfWQolCgErf1s95qYpESrGVFPox7RXKBek/p7lOcdER0/WH6Qm3LZFdn8
F83DC7h9at0ZOqn5Tz9WidH4l+2VOzoSSX/HDVr/XHWkhWQmlf85hox6nFYrOVIVkCRyx0QWLyGC
IBNj17goSPMchBuANmxc6m2LzjeVgKrQByaPggsmiVtwe8ktNtg6Wt8xsgPB7m/htEihKnSv9N4o
d/Zn5ur7P8/TrsRScwKr9qPQc23LLz87CJfg6ET85zQ7THaKibfjzYpQI4sRB8e494a5Oa/BHL4J
nrFkrA3mmGw3dUGfEh3tlrOv1MXbDqIbkLdz7fgcQM8OD4aqMjM63xhwt/7oFQgRyRL4S3KOkJkF
X7tc37D7DqwCYO5xdW9Wx28NZsG1j1HirnsQ88bzO7Wh5Ahd5lZu/MuqJ7FurJ7RAQk0sXWj9hU5
6KFIXLmCUTz5R2l1o0HL6VoaxXrG53PZRjmHaHMMdEWZgqqKe6o3tBEmuKRnhySy9i8UvdSCADKj
fw20gqEn/J0vFHzBpgUFKppkoUw+wVd6hEjKTMNNVPXkMwcTnNizHANjnlkLutLrvIaEFxJElQz6
sFmKAJj1CXiuGL+HejkOdbWlyjTFbl3D1MB/OIvHRmR2TaU+xxR8iRVvyNAMq1vz4tEGJ04t9Nd1
ZWLru5Q9dWsLVoYbzbnM2rdWRvRQF/PbVQ9O6Y8VL+qjWW7lsCZEf0qFxU06o9bYXP1xnDkkE+b+
fLgK8Es3bxX3fEkTkPelMlSIUVeSfGiB0H2xIumbxFvN4dzp3GxzAj44BJGIpjmQ4L0hKspD5bMq
PohPrBN6ish5kH4BD1Rbw0bBFT02awdbWmeMJITuh5wcLoDF2zfgP93OjmsMZpO+zPctTbhYVPaZ
QfRf+FBwjpEhXDOTYaYO2zOagw8v3TLMog0itR8kfoHpvILdbXlOapfO2PAm+AFkE1PMjTgEXTP4
HBJyIx4+kJX/fevn5N7LMwx+6D9i6swJqnrwHcXvTCwSDbkpDwkBoVDveDYbg5DQcjE/HwVEKFK5
BZuMWnj6Jvse3N1+xVU0sRPnTDbVSh/7ubdmRk5iHxFpxKsDPEuSmkTw3/6WX3IESYCApZ/gcxf+
qOLhRBTqFFsiqNEdtRcekrtRt3vKLji4ZfV6vDVEDHqNMF1ntCewHBsurAIhREIpbFl+s1XCvCF4
9mTfWuDpU40HVzC42AEnUcEafmv5KpZzCxrkvFfoW3McBwdUcFHduduYQQWviABHHNUXhl4ezHYw
LmSEmYThsQzcrNmaDB9Il4Eny2RWEuHrvhy3FmA+joPklsOZT9j3prGmgn6piUztaOrv3jkeuM1f
owE2LwEwLiP8sATP3QoiWVHerx7zOJeCYliKxJiKz+kgBdDgAO9HDDKJIEzIafGX9Xm0EodGiCOh
n+NtAJ6aG9FYwsj+1mZppPXbbtkB193o1HmVKuyNqkojgOmofgM1rA8QKFHxPew3K9Fjxdtn7FnJ
Jh3hTU65kdLJsPwCRpIFc68PNQe2UWXgtmtYtON1gugCPR0S6F3ugm6KQP+bsE/v/h3clYqhiS1d
kdAjjTcT+iYnTv63+jMpV3SBALYGZKpBbHfLbpJzC9g/m6TMsIjWgA4rV3lWjFac6qYoqMAt/qPZ
AocZEF9MEa2IYRX/KpPVX2GVL+9azSqO07KfC9yQcTEAAxrZ/p5q1lxx3p9H9Lk10XACTZt7SWnT
+z5TWpe1svmaxqNj9FbiWDMnAA6CQzgcoo9PNxlyzRXcyA+Qeb5mc4hAzk0Novv10d1dfqhPJDO4
HYXQGPKTKEtqH0ibBbd2HbodLvtaLstR7MZCTSXEKZ5CalhEHAZXKLHCsBl/biTHg0k3hh3qFdrx
Ey4ItLXh+GxrkElmiMZA3ocTuUKZefMklIjM427QUGQ28F5Md0dCnWq17GEM8DkjY0rC2f0GZMgO
WeLu3IOs9vaWArUCePraoHRNvxrLCrSCZ16/t3AGqvDD9imCvXM6GCz9jbZxqNHvC5YrnRIj3O0m
bIVLUqOu5PtP5AQmSgsMCIHf7bDqiCdjO4vEnBly5pveg5tkznRJ2LMsxNV7nMbAlyeq/n7Slttm
jWa42PXJAEJClSMHcWj4aEDVavmjT49AXvpPK2BJN1LtF9Y+E3lymRLz3QtDXxamOM8I1jcy2T8K
gz0Fb0biloh5LLdrzg6fTNJ7NkGSjE8xRWxTCk8uaBafiI32/Ok7xKi0zrNapX8OSN/shNSmnQ+C
ZL6Esg3RC2xxVqaqUCdX6YBlc2i7Bkhft6XzlXKPP5eN1q5mgLoS8CRTm8aDpSE2/N34H+1mgiXX
EJtOr/MYh6vSKteLCoNFSvoKUL9AytqbGpluAma4wXZnfd+/jbXZyPXEEGhl93Ox9kLkOo1ss+Om
x1P4tSLPv1cTWQlL2XiDUJxSWGA9jJbPO9Nv9SoVdwEA/VZMdxt47ALDA6KXk7iwaoQLjpMtV3So
XC8y7TZYTdgtNuWknTTWOCg91v4UdtMRtsBURmLELOxfVA00igipt0+bWrQ78DvEH0F/I7LDlat3
aizdC92uhfoatll3fAGzAGvJA4XUOgRW5H9KbbBy3ltjZ9jlpW6i5nPbL26WV29alH1pxbghRcqh
CPgHQuAJqu/cJXZsSIHGNMMlNuSHNIv+K+fvLWFCU5OMXTFPAr9uQxejwadjiKy9EdbTUEOFsdpY
Gy27APrRj6jOeimzM/4jd+OsiYRgVF38ng/C3Gjo3fR5tfysPlSDPireTY8NS5+49r4jFCx4g5/q
eIUZrl2XtIynBFnwdq2QUsIasRgvHKUVCCEB25bzkUzEn1qiz9UJEJsEyoWGKya+mTGSsxJ/K+4S
Far8EbrLGNPkPPtQSLchWvbbZKFKh09n/TxD1q9zXFv8FYKKzdIgCO3RMvhSTOKYXn118Z/MrfWd
bNHQv08R94TadxBbDGSdq33rTqYLhNAN9DpTg70KimJfFDDQwMXPnXVuqdIzDuAAe+y+nO3I//Tn
zYuWwqKTage+63h+3xwnR0Ois9nlc4myq6+DrRVRjs8T8AOod4Uruwd6IyH+moDOnGhO3mTPMHxc
JQtJ6HN2bZxQUKqMXm3wloUCX2emxlFNFojJMJCy0FJiQrIwTa4qZNCHZWirBYteC4iTDUQ8XpGG
JlMvKs+EJlybFOoZNYmceI/luG4f2Wk6MAOdxdS5SkM6RUP8qds87Mrk38Wl8nkVYW1WE7TK7vfD
P5bzdHAmHHMTB7gqyIdWLP0ecfBJqY/axYYlULVhqTnf8dqiLsy9pd0ysSnlnlJ5jn2L7L3ryZLa
JHdrFK9aPMuPLxwh4jOOnYxEYU1/JDjaL0N/GYsVuzS1i4cPTYtv1EIj2NZHGFl+zsrVWryzQdrG
QRblgdSGplW+vem4hPp2NXFHKk7PpanRB/sp2FcwwlvkeHnLCFEqnuVitNmExZ12u7jnvLCB71UA
jVNJLVisJ8Ay9N8gU1FL5QHllw2CxeFyNVdRFvV2EXmpjS2EAiWtpdK2RRK29ZHYuD5awOrtW1yQ
k4rPycaxeruP/XWDjjHvJNoEMWcEy/ymKFLA88ndpLy54tTQEtRcbWh24rrzFgIqSt6pzmm9WYd5
KEc5vCnpBNnm4lfLRfLAQmBhm2mhi9pes42pDkxk/v2GS4pUwA+tTm1Mjp30U96RBpIPch/xX70t
z/yH13O8XtJNOp+W1YHPN1r3ABTV53EsufFFgwD4F/LawdPzX4SXDWfjhz4HOABSnSrpAY9lPFE1
Zk+byiE6gka4v6Fpu4IBBF0MEElR1NuADWi/Zi1+m8mvISVhH2fr4Kd1jq3e56CSqJOoPlDeHWnv
+xS0yX0O20BZRkl4OQnMN3tnYuekIQpjL3uTJIq+UH49YNj1mSCY0+QDjsSvFpmTuwnBsq9dNXgE
MIIAFScgbCWhkSs79NTJcxBWTDuLC6LER9/TmjkI5lydkc9zK4SlGeR/Zz+vJDrf8gPy+On38kTM
zGzC7y184Hv2Hcl2Pgr0nXLf0w+f09lgXniFYjBLu3qeH1yNcJl0DvlIy9rjh1gR413gOIOHXD7s
hTJwfhNoMvWRePHZk983rgu/7QLBH3mwSzQ39o79V9WUQ5bsYOl4dfECQ/sASKeyhAgmMBi0W4GP
myrVdeBzqj61SqKRooDX/ZT0Y2anvgp7hqFMv35MhAx/22tBVgpJtMC3N/36IMY8h0Cglcd82hg/
vc3hWdE96xBXubuxy70zezmQr8nkKgPiI+/o7RguOiSDxc9JTysgvQsaXmBLdcUK0JyTowgZrCfW
vvYMOyHOerX4Jmm+usgWdXg3Lv4zM3RS/+wD00kHXQSgi343IYIHwDyjC8nAxWuw4skx7SB5zLlh
cW3BRwcP4n4cFhc+zxTmCpTQmIyV5vzKZQvjEgEXx/fEZmyz+4eWBF1Em8c2DqYBKp5Xu683JBUV
LHsZZHfZyfV76eUNcM/H/1bQTNYSKQ/fqIPr/OM28k18BoPvJNoEKA4KTAKai6x9GNFTyvtP3kR3
NXuk15dED8+kXHzfhdcheaJrIswk3PUOQPb318HkJ9T5JJZswvB/Cuqb2x3vfpZc2RI2t0QaqCru
wa38OISGapT2II1uUWLDa6vi2lAImS07qCrIrDybHUU8jzvFm1rBzYtuXvj4p+XY+PoR79qI9+3N
2EBjThoa7H1MmEGvD7AxBomwYOu+FWJ0jy2myp+FvlTYA2XUUEoGB0RAXrOJ/u7exbKvYl4qgvCh
3cpBKAsSSzq1qL+Vkr3KUO+1MEwxyNNiLD4GMUfj+gd+quqNqPnJ52/gxrTmZ6j7t3MQsdUo61sq
3hion2iuobbpWGwzHen8j98yjfznxKwlunKZ7VvYSDF9WOLXviLQBy0l2bX10OdnzyHqisbG5PZr
HvIDv3XQsPCqQ7TEM3T7LHWLj3DTYbDuVuGEo+DAbN4r+qpU7XMfJu0l+C6FTWJGLllh3NQYCgAw
VGjbRDTQDHlfmcMjmyvZlcFqjPm689Ebi5nRPbbPCPVhgK3Cd0MurqLlgjgTnRUsD1g8g9Etfw09
Ef0bfKuPbOanq13mrIlLMZZXT5fk2+2eMRq6w57nL0Z71HMS7Ado7Ishyr0e3ajvX2lQmyYHmq29
R3vs87Ga0Q+K5q//nyzrMdpNWerbrBC7Es7qj6sp63ODsR8mnSrRYYtccuRhpZIh6ZqyoT0/jE8T
MxDmyLovI2rL52b/YRcyVmlPIWey5zDfv6pJrQdSbRE0W2ZXHL/phfoLYHUgk/ysSJ7XhINqqYyE
MCywSlj+jznGCAbiJrb6JN/BhGOrqvPk2dvt6xbXWpxRqQRuXx0KmLWESIJNNd70bibYroDIwgxF
sxZp/sq4SOTt/EtKpqmCY5bfRWP59betZA7jjgk27n1qLRNASMMznZgvWVQRc21wDf763p3UUeMk
cJE3EhGi5chTNanI0d2jE4/F5yFDGRpcZOz7J6wlMIJccJlisTRVdK/3xGY2p7ynUzes83MUQSDT
PzhU0CUY808CN24rXANErUmK0Zf6LFKai6kUEmQshQbKaWaPVtMFLzUZYWNIha9LS3muH/XvObEt
fU8WOoCUqMnZ6yYxx/cs6VA4wFb6gc/z6TxkJH+SUStFnSfWxWLesitU3+Lg6jT1p5nD1JVIXjog
xJi6e2v951+SvJRLUMHUfriPtbtVUNhSdwZYVBH2QKnCMtjNW/BZAmQEaLizrMLn/3V5F3hlfukb
F9MubBSyUVYWOXY9BK+jRRIEXi0/2AIxEEs0UEjqW2nwFBSPjFVrWgYWWt4hSU/P9NVyCH9/1uoh
khUL1wwi1W4CYq7wi/5A6uOyp1EtP1kpNiDPaZHRJn5MQmx8eQnywejZmoyfPRS9+oA/mHPPxDhS
x/DtUg6/+vuK++9soQSMsPssO9kSvXrUvWfk1hGacKL/43xbEEBORZIqO2HphVd7GY8FRmkArnZk
PNUapDCSGfx4Fz+wDUKd1J6UvRHmexQolNkGz496UrOJlygV350gseiLkBLr872uWsrU+TKS2opv
/z8sFhU3ky4McJ96CMbNe7B3HVXCRAh6qfxxZvSvvLTDVeAjDEgfCO3IV9lyR0AxyxK2HIehsl2F
V4UX/wIxZz7af9znTmdwO9XwwIY0Sh8zv+JGFUhrSJO+Q41UhU7ws5DAQybdV5tBgT53bgXLK9Ax
98fJeotBUZunOfO7GSwcm6Y/T/oXAVf/IBM26+j6pPIy3sY0bLJhfJNqP2Z4UeBZwyzs1Cxd3r7m
wUNmZ/ck9poCJ3n/4F1P980J4Y0UGSDLgVMLY633qZoS4W/pf3Xr4BU9fNGzcgdgfaC2X1QheHPL
fGtixPM6MSAbW7lFKg+jYhG1wbzVMtySdLIM1XsMP9IloYRpS5MepTFeSZh1SBdZkTTSp6ppIxtL
lF5irG4TAuW7TC8YFKyMpKiH43eNfERcMiJHlMFPeIrcAlrPuRc5VKx8mZaPLoOZuhUlQ6XaDAvx
0Cm9eWfTNTseMuscUeIEAfGXJNFusM4D7P3gAnNy8G5+DTtvMKnq4HiX3RXAJK3AkcoMStYIiMgx
DsVqcH1BJ4S3FGuvAToZk3W16baks4IxHOjEhbtBfXgErpcN3ey/YjKFZMzOXbHazn2gzh8tOhSa
0Cl91OehKoUxpjSDPc3VRsK1fQChLoDeHHVzyNX1PwJAoMxGI4zQMegddabg4x55JzO/xDs13NJk
NXq31QNXW95R75WBxoQh3ztYB2R3i5ApsepxXiJnshDlE0Q2rls0f0wfVqrmMORHrOSR5KckPq/f
/aLyi5qKt8DO4AIBfTw1gMM2Ehe2487qktrgMlyOWS+zbUzUVuf5HeuA0/g9spG/rgi4pNDsrsyB
M8jisunK1WNh1wT6JG2MJT+jj+t+SSrucvQqUGL0VJle0neT2wvLFLq3QS2o4iMYKn8K8ikU/OEh
9NzlYaP8TuRlIIHjWJAvDhJXLJX/KL2bipRqyBdFYUXak5LYMKdZ/EyDKOohwe94HlT2OW5nyI7u
NC4aElBW348TaUnE2tffxAkG9aWng4+y0n7NMETIgUQ8ysTIxp/+d9iIE6ma5LZ8V4jnY4pofWCr
xQ0kmclt0DoXefV9Ny/sHyAcy9ohwwHC0sfBCQdFD3mtNcEZUV73iFsf8CeZApQp2HfKzTwKTerO
BqwQvh1Fe/zPVwNdVqAt0f1h4pldNwO74M2cH1ZJKUtov1heQ6uoS1vfxFeQHSnF7XHCWQkyemn1
ajKWLQUg+0w2mNt0wlrUNR0JTrLivGBN805/vKvb0+215ezbV3JsZuRxmSVXxlw/cqB6PHm1agJX
ESftBoGVWUL+3GFWxSJoeCeJGbjK1IqCEBBAMJmtBEGE6bNYcOB8HXsS56iPwndfuUhPr3RMfHYf
lhSxlfKzHfBro15OQGxhvbc0rFn1VHlseTKAKUzq2L3knXQVdWf3YLGVMxR+yrqY94fa+pe/d3G5
Ek7w8EqDCO9qLqODPYih9Q5ntKJ7LucLVMr6C6gWq9RtVgIRF1RvV2mRZZFR9XBcCBZ8edqxhx18
9Wpxxsj7zDWOA3wFUwWlXSoKauNhXa9M9zr6w3ASYB8H5KK8yF5s5PWxBq87UdTQ51OAfwFmD8F5
DyBBlBJS6a1efpDKu9UTOD85fOUg/2wSwi8D/rcrlgcYqWBh5yEkq+kgpLdyV9ajRS/FKTKOKm/i
9j0lxs2eULNx7DvvqU0OK4Cw4gCRrl9tveDiJNqEQVIX+Jk5cJHToYbwgCYp9teBoMJedli/I8Ol
EaqVzFdqQZeGaTvTA7YqfLehd4QRJ99dHa21cEigdPnDi3mQKFDzIyuPUw597iaaxWHU65MAaV4y
muPdsJT2jSxtuqdgASmblpnFavTdT/C2uM62Kb7D886H+NkBY99RP906l7nNxAj3lFhkpCe+yORM
v/uAJ9rkeoJEsX3Z31610d5fGpiwHgwkU3ZL6HSj88DuS9j+YxZSvu4LIue0JjqEsUHtHS36nIdI
85I93px+TjX3AoC3sNudCY8bzgHqvuKC3bG2Nd54a/R5230wevS2O1NuVkaddKY4IynbQ1r7Jt9R
04WsczhCbX5wJwRCxzNFIzlaor7rC9ht0G8CmYTvkHrSZMrze7qyIXw/uG3xaEX9JLy/NlzXpd5C
wy1l/Ib4EPDTidmlUUxOxAjtRjezBBlXGkCcYrNof6zlv+/CE4FPX63t33cLj1OpN1q6+WAUF4lD
dNJ0tSmDPjJlEISbqFKqzfbNSGHF5KFwN5jYhpCIRBJVK118+VF0tfdKvUCKqQCGy3V/xqQa3fMO
gClu6grPBQldI3mK8nE+ts4Zpi+jOrQpVXa/Ih61XXuyKimZhmEZkjynE83ONeNBpMUPGf7R9+WG
MYZ7899ic+XkHVOqDyK6pdihGNpRiHyIMa//Pdgl8JEgbUpX6U+gwLJFtCaOG06chyv+yeAxwc+C
EMPzl0cixZaIQDJdNsbjCsl0oAPM54KmFpDBFRmLoHR1Pphx+CTSePoNkleKcKaqD3e4M5g2N2Nr
5lZvcXZSqkPe4fDB1PG4gT0sxtXiGezUUYzohRtJGT4pjlX3iai699f7hGHDE5g2pyyTxoTQirI6
yCR65DADwrh0P2KBjo/T1eaCTAklSzfMseG2Xnlw/0j01HLqm/APAit3Wkzb449jTPfNJM5w98yl
ZzUIEqfwjluwpAmYEg8EM5wT497NXwds/rPSlDjjtBMStJV+p5ByJTXDDXtlnzPiXeUfJdVIfU+E
zpf6O2pECmps9Z9swKYf9VqZh4+pfXvqIJ2/juhL+T/2fzSajJMhSXO55dTJoJiuKIxmrdy+k9Xf
LhgInSBpdmMMEeZzfxrIxVYaL0m/uO4O2fGiXxCPfN2J9diOb9z5xYvUqBAr5kTWZ5nnu+0xFZM7
sG803JgSQEOK5v+oJ9yCMIcHOTp9rri1BwsqSvk7X/L2QHUdg6KoDmNHResv8ReLDMo0rZ6EoybQ
+55HRtkgpAX5XXCujXvy4rtGHzQE6EIhntAX9304NkLL/g05w0udBJ8Tqz277CmYehrmk/kjP+tZ
qHaLpiL1QK+iABwS89THwoRX9uwfugYIrRmt5Nm7Ug8c/QZn58/18Q13tDhCIIQ1t+tt89FmGVgi
3/oXTGrVCRHg5SBWgYT9P/oDmN1QntWmdbDQaqEYMYET+WTS/q3WX8dCrsojuW1yogPpIcpb5bKx
8gJpo8Twu9m2oXCWiJhwBYn2Vq1g3IqzxxsdxUrFq5TGmQJIeYXet1a93KwMCa7ywjkMVBxxuMR/
D/w4l83VzS/tt/b0FrcBj5H4PGTlgSR7BPLuOeKdMh5hynuQl/yJBdquP0tPf/DFzF3fEmiwx85b
ArR7nKrasor8Pz8Ih8j085Z1iOZ1WwpwdB8Unq/jxiY6kG1X9bRGfbviPyTJqKph1THh4T4NqiCb
kr8mysDNmXQ8Es+2xLXC6OAeHI1eLlkcFBwJg6tggsOv968+AVavcqLtubWNQgIhVgcvkk5XSeaR
vb3mJdNGmZZSfPSeWgWiFKdiTcA6L0UwlkIyV+Y6+DRkwZ96DUbcwnwmCatH33dRAN4Ens7fxdMw
CN2WAh1dn4fnKvm8NtlBnlpFJG5+/VmjuhrnCGgoJTvYwSas5hvBNkV1hxhUy105fvGee+0+6tur
glLrsFHTGg55uaGDbia2oxht3Ccq5wQcXIeI26JrdRh0zJFGR/J0Cp9dmQL1nFSKYE/26HlLXfAO
mw1jiTanmQKdkWUTScX3ed+yKpAaJqdnj0K3RhBAtNBFO7zlsp0mPRlxAtVplNLE1hLC3BjeSTkI
g3RfKd9VXFQCICT1Inil8/YtQt8ZC1ssdg6F2Mu1NMAMu1S08f7zEEYP8a8efeguLghzXksGoUx6
d7iKTw7OxCuV0JYCshhKa/tASicZYwJjL4MHqYfi8p2uyAbwc3h68P+4Wa+sR648k0xMejRy1njS
RXvxEqoQujf4MZ7ttLnOBAbExPaN37vSo0q6Cr7zARXlf31pJXe4ukCSrP7zU6k5ZT1QJ3iN7Axn
d3PZoh4Jw01ECKQ1TJKSUYZn8DZTLtfEgaKELQQzgBm/CIpdSeXzi57WF94MFsv17pnLxVb/Gwh7
DFuTuXbU3/CBi3a3NbJRTuqIgxPdw9QwSkXZou2ClDbeYNK6ZmJVfZyB+jiAC2h/XpE2yyxaJiph
RhBBmFRjc3OoR4hat2eh5epqwcgw7te/EAlUUvHSjodDygyKc8sqYyycDkF5595KgwPZEkyS49nA
ZZzGmFEOTCID6Zxmf2jlz5u54im4Knn8FeAbKzL4JfALpC4J1n5fDg13asxxKDgz11zD1Fa8Lwmr
uCSFSRQmLiKytJryAbuWhFie/ZJLk3BcH2blfuw0QGpp/l01WzwBWtOmzpmPTn+JGlcSRXMFstke
TbxKWUJ9lWO7TH6BjzzQqERXm+gCyLHTtW2HNVE70DB7LRwLxFvsAaQqkXYnEngX7O5tt9HhJ3wL
ZaQmjjDwYrYPHqylmSQjLqAou4mW+fft/iZeefX0G60HC4dc7SJVTP7/exoximbM5ZFwDHU/ImGZ
ST6zrwBTlDZ/WsLXphPBb5WaYAZOjrhRzs+lux1whFfA++b/zwt9cJEx+0zDYGAMdHK6s/wV8AUI
eoXBALXBBQm45VhHVLCyVUnamaAx93ac7OMRY8khDoxn3VXrwbrBXZ7X0m5uFehrNiTop+y3K22O
sNcWq0S0THVM3CA+6iGQHS2ZkqIIlstYn9Sxu9doACBgaabzQDtiUZFdRcaojs6AkIDUr31MMWVi
ijLvnyIJl9LlLmAH+lEHdCxRHvX3jKMjF8NggxVC/0Uoaf6u64X6+8H0MITBmyXiD705+2jOK+al
u+ZA5YzC6svyUZkT/a7mrE7DRTmWQM4aI0+2ABg9e54qqVerPkWhmVsW1t3RIUojEDuJbWOrLzEy
HMpnJfpFIf/FOUvlEzqpsQaVcM1dlS4+olEKDCcEKv6KdXJZQwmZdNpynsm0vqJqtXdCw9GTcabD
zIUNzt8R2lmAvUzZOwReI/bn4OW44YSeyYCBa5OEL1eTilMR1jpOBcRNm/vCQb4yF8SNQl+v7UtI
cho4CbbHoLC5B8dErXRpWHcQvOb6EDQw9Vw1Sw5ACtWuiuQ5vezSdFqBS+fFQjmxBsBiaBiYp14j
RCoC0Sm4uFs05SmLtxlESqJgzleitoVV3vFF4B++wzbosC3i7UGDLu5AqeQOD7YC65icnEHZK8p+
K+IJccXUNlBW2s1jFyIWOC7jjnqHUhZE/ERXZv605XvMg0/vY2u30p0Dwri2yKyCVreAupTGe1mI
6Ff8Tga91tJb8g0WXpf3MIoOGbxuahxdBG1wocMozcEPo/h0bL3KkF5ynG2qJiM0QHMioPNpvKfG
Xo0zsUH2iVJwJvQ1ZS9SSOUIzwqeiDj16ALeWoMkSAK+2ih/yx7Wzw2+JHerjkPUghwHEuMU0Mqk
EtN+iw7p1w5zx3j+mP1+kmxzK52kCrpkIkB9YENglFnn5PinN5Wc0LOWLh8jv50uDfoyCi7zP3Dz
/ABtj4bgmo/05hWcwdZRPQdxQKVRLWt2k61FgyKI5ENVzcDTZVik/VRZSP8Twos0ZydckXp+kA+K
1ZhtRDXi+ESoFfBXqqXy4Ze4JzmeLE0yTtZsDCK+zZI+VIfVAhTTMi9SLtKTHNljpS3GrxYKkuUF
xnLcz0/BRhfsGBnqDJYEfiS+4fG5tsQBf55rhDAP/t5IdGrdhgjlmRdhm9NGWT3NojVeH4iW7xe1
D1t4S0j/31UaLNUK/hWeiEsG0Uvg8lkyeOvu0iBb25mQNV0ghUxeiYk+EMJDt3AW3FLyQholb9GG
lSKrdc5v18aOBAohQ7FEaUSKYU2WlgH+mpgudU0iROJa1I821IyI5CIpka+HuBJX5d+Ybvnijkze
vlqM7vzTNEFScq9lTgL6eqO9v3k8oBdhA276vzW5jGdX1AhKPTX33Qosp4H7rfgLfGb/xm/Kuw1n
KFDpPmLXOiwuiHT0sCV+PGrKfFPt63wA6EQgtBfTQGWWX0c6f6fQuiYTrRoBRK36WItj9QpaP4c8
ge3uJ7+LbEamrZJwaokDNiLAkal443J+ju7J6qi3sP/YGbV9/okFBO7myWAgDv7L1SBbftTYUZS4
9OuSAbw73WZmZGTTdmgsS0lhn9xA0yI9BoLD5AfrBvKul3rcx3SyQDbO9+DsAJrrJKh3yF7KxdLp
zGnu5YT7HhfK/OBj2HkfUsgAJ5P2AjykdY24881F7H3+Y+xNgay9pwIX3+3pyLUqS0yFUNRIjzK0
yxkqrWi2n0i4tsp8AAJGphqQzwFIjn1zEmHz1pEiVwZizAgezA8nJmdLoT8FqYEtjPTBW1ikEZhH
9iJ4YfdhtgOOlHlk60jdkvx+dzrnU6z18MMvIAeqow58h1GXO3m7Nh7+6fTAQBydCHc6DqVN99Mr
cKlWiM0rH5E4FkAxkperbRBMhK+3fvCk5jdtJ3ViUdZdMjjV8RlzoK/gpEZc2mht/3PubcnM8Cmb
gqrBItVIQMmkfhAgD5ybdv48m6k7+6uhTR0qiMjtsfSiQpcZdPx7KB1RbdqXmDWC6UMHIqyFR3m9
xV1shO+e85Hx9a8qwxtPBQ4sLRgn9LKWBFNzNe631y2uzdrUmd8jNTXa3b7SRAHqZxTDkUUXpyDI
sZBfQakhV0hevKImaxm5cBsuT+yiaUg0wZ0MVGbbcqcsOCVzpYCpiJRh/FopaCpZFbJMWTiRxt6s
xdbfMLBYetiYBJD6mZFddC2CKPV7rrasRv2ngh0eZx95SID8GDDwg6DWubUhIcgrSBPAybov7+CT
P1SKmlkifymuDdOS3g2XfKAmMDPzZqmKQhfS8SphN7EIZ4PKawt92ssZ8R+41py9w8UzkWdzuko0
m73JFg9ajO1KubLeB+ty+3hLbeybDme7DuMfhQKxjJNh271CFA694XAam8MbFEC1T8EKYbOmMxw4
jCMfk3+XP3aYl6wn1UVOTfeSilOyExDz/eiTr0eoAy+MXU0DlgbN21lE/m8OnMcRE6f1P83ai8MK
LY+FlKvjcIKKlKWbmehkBgjJrT2q9ZFIxyfXr4x3xeL8IKD8YXhE6ZoyXOPNsp4J3mI6LLHxIYMv
0rGSNhNQ6qMVfukWfYU1iLK1bNbehiCoWXRX4mWmCI1iC2+Y/M+/x/QOBpR+D7AlAi4F+RcCPf1l
OypH5lpguLOFjc+Ej9divBZ6MUyGx536H3+IDylI45pVzdAKp7RqnjrXt8LhNt4iFFTz4xoWtLeh
c0TZUvMhUKKpw0NoPYoD9OjVt5cxxwxLAI740+Y2bhlHK3mGKsCB4i3wQ8jJkvhf/LQKKl9qkGQ/
NoYJso8vOt00R6aIafxRFsWT7609iHENanZ4Z8Kjz9sf14biUWzfcNVKoBj397h80jRswuCyNIKC
dDDaH6YkjxdADWBCB5j6RF2OvnH8LOT4yQocnu3Zg+OtxD1oWQMz7kyF+aO27zQGrPPSoN1rF8G7
jGDD4X4zCp8+FsjyXdqJV3n8hd6gBLldbLOWQpB3uelhfhcfVjf27iWGYxlX+51UQ5igh3KkJPUy
feHb/Zr/pYQ6XI7xc7ewjzAJVa2RQ1ReQEjUpzgNGRmcZKKhsp5DDcTCYOsgonxZVmLV6stUV5F2
PyxufI5QoZTHi7+dn2RqrolNQ6z49fzP/a5quG9hnD3pz/etX5fdVB7uJ1NL9aD24wdFCECxM6N3
Ky7NqBxR+u38cBFS3NTzVBY4kFSOy3ESqbrmQ5/ylk18tbdvhQiT4KZBE0REpUU8/Gd6a2S/1dF9
qhhN0j6kKN7jgJDQ4i/M1rU2F3R9UCJwHU9MiGjBPdTDeW4MrPOzu1AHXe50aLdHdR5gtHZj4B6g
52ggAmU5OvuA6xI2DnaCMvykVSvp3f5ygik8lcvkKsZHfCorQoCRVoc3T7jcukGZD9pGWbmsVJ9x
sFSHSz0G3ov0v2PnSa2BxNhuidZ7GtZui1/zVSKD6pM52CwvQgtdKW8YlGYBSVFCTtY2LBpRjds4
Bfs9/xmWTtmTASl//ZuqBW5iThZhfbtGP7M9A9HbWZZqE8ULYrybUvGepOrErrDHe2weqlK5pAQT
PQThE9cS+vzLlvABq+jvHsMlu25l0isnFgpZRYxIg4q00aOtzbVGHumDgSLtr/SeWC6/tIJCKPhZ
rv4U1uNVf/NYzQn8y42x0Ldybe6Vqy5N4ZjJiMbdKXrReJq1ZS5Svkzx+fOocSvTreQQp/YtQYG9
I/vxATo03QMAxNRAvcgeAo8LoSeCEXStf6faF8vZ5TxPFdiAuB+DvX1c2sk4FO2iXPPUNgd1Z8v3
2AbmyyAUBliGUa3W2C7HVg14pg253s2/qmCU+V97cFPFAAhPqD9G3ckruI+FXj7FC4+IBuBPo3tt
I096Gzbg7pUDglyWrjjno44GxGAbaz8//B0Of5SZXADqnLhI2yWuJTvmkhsKxWqG9LIlgpkdnNH7
lzL87K0JDb8LRHeRYzcPbhqQyrWxs67OR21lUx2nvfd5K0xO2M/V8hdM0ryjJGQtGFuzYHBrNXQd
XxeyHYDw9+LQJoBTG3IgthQaVMC0jITmpy15EVfKVfnuy9SaABaUueJgh9mEzocxMa2PPkNZcKZD
FykHF2m7EZknhenM9SsjmQBuKJGyojs3LayAQoJZ/N57sxlWaj3v24/aN5O5wqzezPfnRKgLWaKZ
eAo9CxjNHa1v34UIwB6scxLJ7RDGHp/K/aVQSPDOAEnTB7lxoNa+5vMNgOo/Qo4eE1hYN9AlZknY
6IB2yNr3JT47HgschCDBmto1IB5xgzHeG/WbpE/lRn+EqzxRFrfae2qNa7+KwUeQPVVK67OpQ04w
LZTPL7d2T83xTCtVJzcztMwLGgj4N2/N40zz89HR3hjUccyW23VA3RNFfuJB+L46Tz9K/34cwcz3
J7ZcDFQsK57HRJxyKwDyWHc26YiCHRWJzTG5U+Da9cDwsT6E53Jk85yn2Bc07zVBV88k9GfCd+wg
tT104lW9SBpVTpcgOvVjvG2g9YGoEX3xlf70WdtfLrxb/GFGQMZRfENbyv+M+AjUpLvrYY43BZlE
4Z9KJ7dGCdGyjBrC0DkxrsHd5em0mDiP/W7hhSyKRaZmzi8Hsnofy1rLSackYMaodOfRldG7Ckia
W/dhoYGyV6PjyEaNGtCOZ7gv2CabTg5DZJ2c6TgWUmYbFiA8BSRaPgJUUkKVx+PWM0NXbz2zkN8Y
5K+dkYXubMqSqAq0+mFxWBOGqY9Z7utHPEq/GjbNFPQ/JFZjPGUrog5/YJEYDIeP6v83VC+W/vMm
uTBbtSkZQ+O5bXGMw9GdTeLA0Yfj+dA16r3itymMAAi57F5kKa70bjraGbIb9ef05HDCyNMxMnMw
cEPi+mjzJiIxrndipMeKJKpOKRsKn9tyi/3eRxKgNWUaD35pPGoGbs0TOzlMXEFpF2u7G/WBtkrH
8Mi+kJGljRp4TVPtmzyMQLUqRtAb+qWg6bTGVvicINSaY1MZz0PAVCN53Jd1opofcF9rMUxB0L4c
mJXK61TZoXjDlzmpVNut/D2GsMJN/03d05V6QxvZxSpHS2+haZ+qJSTNe6waGTxwLjHF7KNDCgSn
QvkV9m0yVgrpmlkB4T+mN1nKdfIKFNPCmXlVaRX38Pevk4grobqnJ1/eDJAiN2IzmZiIUH34NbPS
j5VG8K3SCcUppn3TsmrGXEO/vxkTaos3lfl74EiWAV7HJkpPM9O3tsH+yGbwDF5cjJfC1nC0sMVg
ctMalj3uvqJwyqXx4A3/lPeFgX7efjgDJIa0gr+ga76XZAyK5CLxwzH5w9kTvgiQZqEUo5JSLFYq
pfTSrIca9cmvPEcdGQ9tzGGQDIOxGjwaox3FtDI3Y2YpJbG543DSWPOOEa0Zcuez4wBnvr4u6kQE
P6JomjGjAHNutqlPmSXzZMj7OmKK7FC5bPx0eIKmbAtbF7p8Q8htf68/DPdrLmoM8irMEaGrZtv+
SjQXEjxz/nIJOwPjk57rGrjC1UbTi1ZS8kEysEheZnohI0/8DaqEqItoVq8xFQVupJ178B0WtVhF
Fb7Wu6nSMUiVhKZST1avJa+/O+1bXQuXpIC6hK1w2+G4a4QYARkdSStUAXV7UwOBwoEugFe88WJA
i/iepI8gyYl7IMGCstL1HD2VGhJaPaNqZSOvrRzSxGB2gBxQJa7f9vg0slmsMzmF1XU4C/jG9tn1
LD+u0MNMo5voludzz+BsyWvEdIJ1sv4DHF6DdgNIxzmUMrZkUOyAJRTFoVpqDqhikFLwvMiJJwcu
L1PToQuhrdeQ6NipUr6IR+wgUu5oEvlmv91QcbZtkpWz1wDr2gBLN4icXLRC7bFdCYWGOivwFcVN
RszImetIWuPkwW/G0xappJnb9BIyhEuKaApHO+LBxYOBj1BAdvQjHfaxrwVkJ1+criC/CDLM+HF7
itSsLhwLQfvbB0k0f1ohDfVSYq05hAbBJiCljLllqY+cgMsVyWTEQ66Qh7EfvhLrYN1HEnLjbfWV
8IP2nq/lil+VQJ4rIX5rbMTLOmu+SmXmVY+pFgAn3jnnKcGjl+v+BGpq1uqcwd3q7zXvXFBsTBu9
ZM9W7xrzcpBEYM9It66TenegsEhXQ8M4q1smi3mtdlD4d1YkOuZ/jce1qSLdhW2a8lo75emuyRzM
U+UlBz9SDbUFPNcclRMx9njDvF5SEmUI9GPdGpcrn98GzKnT7nyXlSVHyJ2iuyhmY8Hf7Uz/ipL/
cthTbEKYbSqBNwnuxcUbNGvPvTABiYOzxN55VNL5FFMDCNl+Y8Oyk2SrvBLmhYns1Ch6/HzOjKOc
LE9WLwwbjYOKYovpmMH4yUu+TVm8au8Y9J8JSvcl2RwSaABgrPX+WELL9KYuicp+8ZQj23Hv+u88
RfZ3fRRD5hkiIUaQoWkKqnZeV28Cj7YZleMbUoU56w9jxMjc7UoLiPmAostK62Sz0rMM9/ZXBVC6
0pHEdWK7GoC8YpcecA//oScoKtujweyC6OvcveD2LsiQ2/bq1Egog+B5+cLKxZg91hLF2Z4OS80N
8OsTIDrEoIdcCgdHE7Cj4YQf5JNkf0Xdxr0Vc8zltjbV5NinsSfTzyjPK/aN+9mjhhtYT07GRbCk
XnQDFXYpVxB8tX6caEnaFhFs7nABFdJi+mAAoXzKbA3GnmJRCy4zgcf08Mr5oMo88dtzN74m/v2p
bzq7qABONPt/+5hbtSy5tIRycG7D/7giJPi2zNI9IZpWNaErhDyv0rHEWupuNvF5X8PXoU2iZOw8
Y4/uCpmAhqgLzr2BAUlr5lvd5VPiCFumyr9PaXnj8FKSjosIhPEeSTf/17G/NKJAkrTeDyE/2keg
UN6jN+efdDgKBmOHrgM0xRIENexMt+z5cIdRvw5x4iIhkloP05NjHYJSJuVK5PRynsnY4QjdEQSj
CYnWsnIYSTaRniZuoUG2hurDBzsXBY7VklDCsdnl20c4QxCtNkvFHxkZmcqq/JiNq96LDnkczQnR
BiC3lHy19tIOPRta1uFbnOz6eUTUtlQChUAM5WdAQ+O/0QJDuUJGkXxaKF30olUq4GujuSlOE7oJ
nbKMwfCBlVck9Ef947xinLd2Tceo+9ymYJTxt5RvuU0KL55GFQYRMJ7YZEgISYKb50SwTbBi3wiw
32YqNUVcpTlr+L5yvNaNOjbAyVGN+ICiJ7cF83uacJLE4DiZWSDIa8CYWzp2lnVbmVv5gPdGDwwx
T4+218c18wGWdmTqhKh5mZAZHp2MOJs7j4Rq1qwqc9HL7AMZRctLEuug7IEOz9NarxiIs69bGpCY
sZqVQpkKUJzY6DNN9KS7XjwgWMa+0rOg0pCnlsQTA3twGFfyhKmfO3CIXt4Xay9Nkf+faqM/R91c
Xv74vZyaif+MgGw8kLB4+zJLpTm3zoYFzluVBrMk9V++jfjijsGEfwzRGJyGJo6b6abKs474DPE5
vRWyFvOxZy7c3N5O8It0jCkGCnxEu94h1KA9Ar8uJRUaUPDngFwgEkJ8KwHHoGybj7niHNzN5ZLQ
Mr5shN7J0HfiH1CLwjV6oDZTqS8GJcgn2dDDR1egY2X8pXdksKtzMMmOsVbnW29xRr0CmVcCVUSI
X09QBAxzFyFXYDymUpq5g4kvMqAQfCvlPAZ0phcbUUl4DuMHFILhkurA32lTNv37f+FkG6KUxKey
NcCtn5xlbX10wdj9ypNxnp+IgML+y6pOyDmUCIZHfz1LGZYKwQhwJZsoO0RbBVIIg7BYKF29RD6V
3tu6KZuRQhu8pSyyPC9CKLeqJe07TfaPmda2u0MYhsQCKsyWlW4WklJnbSZWSBY4ho+ouvr4A+Xl
wHUwbbnaCeKJXYOjRQeA3AS2PNajo2OEJ8cCjP5qKrT9yc76XZllczMlMK3UoST57yVOEfhP8/qb
g5j2YpzeUDXH9qHIICPQyjKGCLD/cci/Ni/k3or/KPpR6Z0FaEkI++/d1N8RCnbQV1dsZba2v18o
EnBEoNgbSRQ/c3QyKNQo76xVdSWV3Hr6+9Owz8vvhzwTL3lf/ALx0Zop8oCGQfr+ShhZH6qjmkIf
Cb14EVR8BE1uRTthWTjaIruse5OwN3Mu5cKTtz0m6xhjxT6EE6nsoWdo2UtTAbjrWMSCSj58fRbM
6TPoeAnizjWZvLOM2Cy+4J/MQ3Z6kvsFr1bw56kUP51K9JmWmWMZ/nDlgapSM1+0DurTHklDF9eX
Cc0HbbKLgwyqtnlH14ZGcSMrfbkKpbZD9Xgn71PBAgZqgin6gFsXA6mxtWWULdEjJX0Z3d6MfXk2
8QbogPjlPx2EXiAkjHqSQPxMSEQYl4eJAbxy6S1+KBzULGFPvUuJAzjX1+W2dXgUXNL8JarGR7oG
KNlTh4jUPUDQkR0nndr/GJV3hvUTLQGd/12T6D4dvVxhRE+yfpQx6DbF4Ej/h6ZWn7ZORSn24V4x
mnkpzVJ7y7WFGY2/Bwuh61MCBm7BxOsknfKsvV1TapaLOKLkWJlIepEM5Z/+5L8ZGSz+ElbTHV+O
4r9aMpCl/+D5Mj/iC32M2zcmXprIq5XOo0w/ZYzmxkFkYAtL8ffhD96/NOVuU+Y2W+gfmzjdKKnq
qgL9E3admELIYuBt+6JTat2zcBswfF7pWY0+nFOnrs8uBzE1mXLqBSHEC8fG0fxN+WuxWgaqZQJU
u7oVF2qUrkKA3S4IWwXqbvQkUbrNL+twmRqkZXpyKNsti57t5vp8EclozER870668yEeh7c4IDA6
nfplalCZEiVWV1jCXg+lUB6YCeTPG0pcqSosVwCisPzSNhEEhWzi6khBW6dFs6/HBeBS1+0yUjFH
dlck8YnYb1WK3HGtLMOZ5w+n+K2uGBYZ1nvYF9OcfR1OQS/n9qiffEF2tec3BLsN6i35zI2LCJhh
lcI+3ZnsrHIUGjNAJr9RD6wRqRfVdHmFbUFNJG5gJk3XVv6yk0FR404gjpgOb7RtdXcIfSqmiqjF
hCB+HOy9Mw3vv0c/HlLM+kV6EhgU5LUKE2C6AGJ6gZ9m7WJHwgYfOfwHsA0AmKbbgQw1RW5oDQWZ
jFH/2DdHOYKM1Rv9m8PBzp4TNijLS+X+FfUzdP5/7UKtQIJUSh033u62q52X9RxAEVWJBPR76QqH
IdLI8Pbv/EYDcIC+wyNajfwwNbAwKpf6bLg4OAKwRJIYTm6faeuikkvIHjZy1bebT1NPawExRmqS
XLJQVe0iOabETtXouNF+zJCn/joLtobNIQqmEAQmMtonNhkLMCSJat51BkToGwLdjVAZ1S8z5RSm
IzXGNUmX/OnAwBmhbDQBWvtVA1XZ3UNtkNove1EC/NQLRCPrl6PI/6tWToPvl2uOGe+dv+0rncH4
WNZ7kSdaRqAVQz3+VAOp8JetPVKHiT5sme9mN4BvgPqfPilJqj6Msz1Mm5a2FzcmL3VCVIyNpOr/
wTdsL7IzRo8c73iWB6kRoNQ3ou4Y5qPCek1alEXoPkW3+gXb4XkjkogJ3NH3yZEgA9rJEHu/TV59
i/DJXiMIdqLLmLVPIR5rkbGr+Bz5tQZyvpCsaGt8LtchWAHTUXJU5jIjVcmwqxdvjeNrZpNxfN65
RNpu8kHG0gxokTTJq+jPXLVZxIotoikPdVzg8yWiUyBpd5LGy5MSrYg6dF1jDkKnHti+rVonC5PC
FWBWr2qmWTrAfAjf0/AX+GQPbPRminlLEVv+O7v6taVtmg7XO6DqEBIn8LQO9PvcwIl5YTJdZZq+
K1Vov7nP+vQnXEwujpPjwUwOFz0egnGk0reLlFZ+HztleikKnfqqLWfwR2XMPY+KvrZ/y0VuBs8f
woD+u0yyqZRdcohSPyJEb21KbaksRZKwFZVVH6w4cKTau/eWCiw1QBoCrLvRD5Wp4BxUhFMs9x4u
058vzIFFn+KJHp/YziK68i+Tc6dsnRJyXc02CMbHWsqNFcMOIPn6BEWanK1lVqGk41hybMXUgK5U
johim9QPGorzLSR/SodF6vU4yoIUq3sQcyACGKonOySin2ybMWGv1U8/n7xZcON9Y0G6bfjmndiM
OqLxxm9S1VDOKjCow0mFkJTXONp23fNUK1C98JBXBK+GGMUnLv6fq9XtIexm4wftbdDS8MJuFKSL
FH8bUmyoSGiN77uOsBs33FHhj7TzkQY8hUybxVfvTq1W0Za8Bbfagocu2Wk4h8inK0dXz41xizQs
sTEHVJ6VuVeuNMuuuyLGaTx2VZMtkRMS/rHTp/0Zti2B4LUuErmunXgt8Tcm7jAZcOhJSC3tuX4L
Xm8jNDH+ZC4vOC2gfZ2nthBQL1dhtxmbJkionqU6ZGPKk45Aif5ySMCcn/Opg1gIjWsJwFlVJAwi
SwKF2mgmOqo1p1FApjUXE+ZhcVF9ALtPHPzUzRuVSSDcINX62hUbvecUWlQZzBBmN7FWfSlzIbdJ
O9OTtaIOawDmMbVv3IbqH0wyvRPRqIAItZV3UkhDILaSfVUGdUanaQDrZtJcHNaYb0G8SJqMYXaV
aZlKp9DW7YIcoRownqfBLTEurfyXewKSvAQqNCGzhzwPO/Gqfx8JPPhAxC+HJ1hwgTxXeN8IbMF1
UBMmTCxysjZ0SKfxdd4jMfB4250A2RajsScuJzPzSoKr7nwIkhRQrL0Qx1We/HweZC9aBzQJ/Ahm
hLLZoPFlKNPbHz83veuhNk6T+V8csreTZGqf6ZfLhnCZojL1bXP97d06fR02JyGpNMoS2rSyhpyW
LPqtGDZKRBdycEaHAKMSSAE2D7km/RZ2ZWkcchVzEK7ceNmGe1rDcKeqeR44a6+1ZVJVsVcyC6jC
0k/Ivv5EX20v4xmDs0Qq0CVYx+/6AzQEsaoAVzIP84QmI34CbVsEgO0z6C3szlMntcgH4hn3H2WA
n3EuHzKWoQU10y9gSyiDEaipOUrjx/Tz62vXIzYDBKEEYp4CS101/hTvyaCfoUhSc9OqEDL/M9P7
wKcmDn1X3ziBg0e9AohI/yJjAFYWeAvyEqXr+VbX1Rh7cS6Em2EZkLNk2wEH/n3KVKwtt7gB9s81
hPZbJYG13gWWOXkSN3kiSzG4iYCi2eHBRvby8wHlN7rrK3FzgXgFMAXB2D6GIeCJK/OGdKBUnEF4
mkIua/gs5j45+FwDt7VmzDyJz4r6srzV812bgm3nqERMqiLIsLcjivm7fwL46tusYyMFzRHcTz3l
hafEkjvJkTav57/wZSBFKrGVam+Q/615aUexwzDV022mVOXruIN+7AXxWf2EqnyJ3TYsxqU+336P
rPyJ1PnUXn3Rhf7BwHn3to0E5s5Hh5YZ3GQzv87kNKWfCpl2l2EUDjeRYdxz/ItIAf9K9B/X4GYF
cgyHjFN1VRNE3RJBVVHA5Z59QLx4ksHP91askkvJ5G5gOZndxV/eN5wCb8B9l2ZGqnipJBUhH4mQ
RQXr8/DFDuvGv/Fjsk6oggVSHUW83vUYvvovaG6EeQ3WSyMU119NqdMhIM+CfrIe5ZuiG5xy3VVd
2T9FbNBBtKZplfS6G9dAg1LGEEON5ARUjx9AIyj0J7gr1iHsFD+MTnx2oh05DjfxaMwvnEkJ+QBS
ntxQ79kR8p/IgiFrZ2AiaMJuBBP8wvvATVTKgYjzTlOJC76gSwaprtpFzRdKoAcjU3JRQU0qbfo/
5D2ffNNhi06iZLrKQzfDdK++VzC4rav/3teiB6K+GttY6ciRQa/7Ey6jJFFulBRE28glrpD0Bi9b
hKisXLs6qRi4IJdKICly6JeKnTmSOqyepsj45zFn8KdieleExg9tSK2fPqjOc7os8QbxQ7pd+zK1
QphR6KbCwZTIpHEPUxT373l4v6f0ibd4xjLXA/1kOhs4ael2aIPqlKTLfQReV+4WFpG2gKQVzLYp
pvaU5zlCDITeVab8QIBEiZqcWEYq7NyciffIjQ5jHzU/lNbpQI5q/IIah0DooLNyBvjxguxa526h
oEXu2dQaLg/tD25hg6MNPYi56nF5fFv+ZEWzdtZ9SwvoV03hmCX3M4nQCbvmtt1zM1d3jjXDxQQH
rBwa4CIhL0NDieZqTlq7SKMfvACgEBgw8PoYWbaOi6TvtkDc917VB4ugV7UbMuUw/6CFawxJERp3
ACQFf8g6eE/lSG4uY6QinBb0aoStk1d7lIdEj+30WfDbHvWMO/0SV/2N6xuoHuGZMMA/zGnLeJsx
ZvuDoyrBuM8dBGjOCdijzWRi/J7+SuJQMEyiiZVRlLCVCo6CbD/ikLo9iqBrojjzbYThRT6xPItc
wgj4jAbccbDCHozB6n67DUiIs4F7rdTSmCdJIf+2mqQsEh/zepaxlF314QEwCRbmqzHjrn+agzzz
fUnybg2J12GFkhsU8e5+2FYLPi7LQyylQDOdCklStXl0TnLav+TVf4LTgcHavgWK6mLpZruF/ssJ
k/L8EiD9pG0EficA5EJNtLdTGPwyzh25HSo7n+mDuXZt2EBjLi0tpGF+TQoVzFF6TUKvQZtQaG/W
WGlg8CqBTUEV1Fam81tBHXI6iPX/IuNr2LBrY7R4rkY5malTNWjcLFsi5e+/2WjvyDTXoUPvHcnY
kMmxB6Y63L2M4WpuSadhPp1GeW1pzBJ4uG4yMBdGMy/vEKPJuUzC+xmjiNO5UB7BUZQNKBG9PtsR
GEbwo+nX7fR5gTp91bXTcRx96B1HUFFzjATKRFlP1X1rBBDH+Vmff3XndbTdqLQDN76bb4woqOpt
AFIQ76R8O70FTHb0JLJhEGPu69YuIKKUrxVsnCjWVsxt8TRLfwe3XMv5fF+h72+YVxE9EEmJ4AL+
cOftEIXnVV0jsEDH4ZvSqaDDGjMRYsoOdLX45WiI71YpwfqMu3PGu8VWpjK6hb03jKlC9gbQfXFX
p3pEzVxgk+QHqi0ccpcj/45OM8vS01K6naSdKWJxA36h79xzQQGOh9oovE3a4Im4KRHJX99nBHG8
ZuC42Mwr2cc0/1o5k64eCcUHmFnMQ5cUVxevPvsHT09a+TKCgUJmyMbqtYU0XGUAslkm4lJ3oAM7
FXDEkQv8UbVYd60AoFbvx4mu7vfHEq6WOUIAhuD0FYGQ/rnUFBKU7uAQVjjMcWjxEXaKSD46i2h6
PciHVrF5rJ6TTdobuenpS4De20UptKytOH75HLZTSyXnh0kC2tloEb4zrqmqutHSsz8jn+eQXfj9
a1XpWAFpBbE1192JA5irb0r7cnO0o5jIbfUWAfpUrPq+H03/Lipgzgly/jc4v0CBUcCkwETf3Ql+
Mhc0u0R6TtXq1NwnfMmAePLYV9lFa7xzS9iv636pDr69vKZ+mWcsgsm5Ki0MVjvGI5d+6Gsffy4S
BB14OVOoRduEqVe71kjof1GUnXg3ZLBVvkeK+uXdd6HvC8rBHTjGH8K39ow5LFLJob/Y4+VxS86K
MHUnRYBGIUx1HJzZey30MuKE11y4k/64pDDvKQm9WtjltqyZ4tOf6OYl+2WEqqN2976/5nW56THD
Q2yxCfjGDiK7eIP9neWmZcRoQ4PZWdYwku/wjoFbq+ogAIj9fz/SB76XSpIbxiIwo+VcyWwet1bP
TyUK51sxOvdg0cGrOm4N26dGlmV1YN27TMc1Vu0aQeQeeqvoh8m/07XEFhrLEwRozF+00xdv52mp
3ft+jx+XFky9PF5nnS0GNP9AnsWYPikXu91Uf3xoa5w/iHTj0fnHjkV6/D6k5y+5kOtR7I2AkFLv
zZ09jfi3L3uDJYuLKT6A1/hSieEytizlh4Tt7U09DNlo86Mn0h4iu0X7uKY7uzSkT33qHXdqYrxb
Wp3VhQpQ16o9wJWeeVQtKwu0jgpUOOiNVwVNwS5wz3IWM/tctopQ2E5H5dOVnjmxnYJMFwvUVQfd
tx/dh8XrzK2sC13XlhDFThR7iV/Kpi+SQ/Qxmj5Gs04JZx0cIdMynsKHeyrRrq3G6pnHL7lpcdNv
nFUz4b5iQIkwMdaFVIJ78TFhfV4WNSTcu+G5yYwvokRRA/OFxPIhKuIANZ9ObJwczRoI95tadkf5
nCLZqwJzeltV1YDPC6vFqJZRGWm/zRnlAUbr89QlVqfrDclcB05J9czTDKHUaMPR/yhJvmA1Lj0w
jETxbAcmt3CW+dsXiFZfLxPPNOXdFY7ckvHLWfxotChgVmNZuYj3rXy+K5WnYBB3nNA5BX/Ky8st
j1scFAHx1vaalyoNBKDHAcafFcsvJ13qk2x2B59+Z5aL9bTujRccp0gmWdUJzbh87OKrN8s7bnY/
Bt6ByTntHH+JtiuFIJRiE9vmWqtZvC4D+Ydtezt5ngl/5v2RGec+1/e9anKZSk4D+8SR6Z7Wum6x
71X3qCEP1MiVJzRScm4O3Rx8uSSCJS+cTkOakjUgYImnXD3NtD7pSX0n0o0Xc8h7+6oA1Com9qaD
UH5lDO3tIBEljFb/CZ9Kwf+4hBxfNUV4has3D2/0ht2wcKUuMmCrK/XTTEuV0uSk2z93361KlsyT
99wFfWVhIkZ6030ka2MvBsXmuNe77nCW194C1nSdP7T2C2zpx1ueJeH4nKn4AYqalCoPiwi7wOu7
pFy+wuzgMZ8lnRHd9Ct+gnffOJ6P8VV/zZTrQm/Yg6cNknaboKfKgjEQD7UNU0EzjDaQbOhIjLq7
AfWNhw8raAtEsbwYajdEZMmQtM220CbNtupvfMWUzgEKdS/g/N9kfKHyTKRo0zDLGk7vD3o8rNMB
DX95ZCeZGGN8KI+au1u0r928KQORO836refkStQD0dopVEqyU4np2JUL649ek4WcuQFU2AyayzvV
Q/MzTLHFBZDYh+S0K6dPcULeIuao85ElIYYY7PIlVNQAF6jEsVWpS7Sdb5N32croP5piZ8hGT1eA
l0rvsjEIN/SKEVoAc5c3G3X/CVa58O41aFVWpWRwehQmCXGsgKL7lRWAjkEoAPw1PzWtQQtZBy1w
14Ny0yU0PlFPrLtYhyYrkkD/dv8+SSKM2C27NSNRrptmDmdBHRJLTYMwqalZcMsOn1GP4f//gPZ+
ruVdoqQ49g10RaV/IvH6G6lvEXxbTKiGhFXJ5umHTnqL1ole1U5Kgg6ydRxQYaw4tPHDsecerDkG
bboBNlW76SoXQY7dVqF0twMLPvfNwTEeCbS9zthX497FtOs+VTRJopCg1yhqXNIW9f6nJEYpz/uV
bVruVPPmVn/lKDR8kemPp9FuAB22TofCFdwljEU5RD0YdyPQHGQlBwBJIwxr4zEehnaOR/wTIu8c
B7zwCIQ941o8vXpWe7naSR6uJzqjlBeglHcWLLQ1zpMn/pwc70pZRzoLfnd+pjsoxoxo2J1nuFeN
rZeYRiWFgYs3zTJLPU3c2Ju0IU3g1K7AMskQqa+YWreDKGUaQvqVn0TrcwtFTuvfFbDW5/qiKiQz
XUHs4EHvpE5fv/5nIFDvVDxzRMR7Z4uh9QkLrzxFrsVbtEbQugDEjGdpsDzPkuUbza5XSLl7/hjU
S196CrTPc/Ij4VcOsGjJcns08M2R/wbwj87uLzAiewyD9JnwOMSETYobC/qZpsHDr1Nqcbh+DrkQ
WiJAmpTyFDSTXF9Aq+KMYt5Xgxo2NslYn2uqpc+OKr6TsrtIzX7IVf4GO2ezX/rEITqdky5ifBwr
o0iC66ff8eaSi5NT8AMY8QX2+WTOdg03VdGYbLpt47NnCvKshrdJZw2djul98+R2tkqt736VDP9t
wZLgbBEfBVuZcAFoHEDYX9ZZXcY2Ad0uYz6DNcovAaDNdw7/IgHey3EQFW08wJ19WJG+IIUS6Dkt
WQtlhmp/kJt+I0OF8I3FX1981POUBpCF/UuWve04kB3kmSnfp7MDe16jPJlttfSG/M+co2Rp9HoB
Et6PeY9xN0Qt84SYFybYfF2POjac9C7ySaaVEWrDR7ZnUehWRazPg2qPJnniyI0p9mniJpEdoRBn
5lKpjBuZkoSGFwQRV/CjdWVw8d6vZLQ7EnS805n7MY0pseKtiu0CLlk0DRmAnJ3W2x+66jCcqii/
uYsf6xTNvDpvEWuN7lP/KVf8KVPP+lKIIq04Pkl8pIosbfav91IgmSUqrd62HGq0bMzx/UUTqyUQ
brMvLoFoJofxNYPS7sO3MWD4oNMGRGw5QE5Ea/lvio9gqQ/i36OvIVIwMxbIQVjwxUYPHY0qJtMX
kfXPKdxKQphgN52xbiBnrsKsmOO3qz8jk0ZtSM1rtl4Y1GqumIWc2/degRB2SaF8Mt7MhlMJectC
1Eh7EzdBRXLDu5zyBi1tBDKRUDE5ZmXcuU3GbdaDftyBB5yIRhd/xrZg/F+aeS305YQxgT8reY+w
EPhehee2z6bVpyybQKs7MkiU3Em/EwMIYE506c8qfgQVyBrB9TaA4Bq7VBnmmf76367mY3cgUWVk
oNeoaKjKTa4mNhdA4R1OfMfXYZZVxH8tL13cjhGhlfrx7+NU1WIONcq0nPo+vgNh4kuAmgwVD+pm
0V0xyrWguz4aaHV94ExL0plhyoeapo2iqJxJawYzo01VhqkZN8uAsTArAkzTbc4telTNzh+9Sd/T
3JO/KLtXoEmWGfElIBn2c5D5TfnadDaMSr1nkw/QAF2sTWAdCKpXArGW96aoLOiXLTIaMC4hutNm
vZT+1Bq/BEd5EZ/QuVgGXSjJ/D4mXGZXk4kdeRcuTOtvD5XEXsPD1ZcWv/3pDC8jaN5vsDgSk5ev
nOz1mFZhyj/ih7enipj/+lO3zZ3U2ql2GD2cv6jNsqqMklFNi5XjV90LMHaeK8p67rFatir2ggku
7zagvtU6wJ0jUsIsj5C0VmhcNpEH1Ui+T8NbWXGcb6Hki8Uk6ixR7YF6WqVynGI2+a2+kDNTA28Y
bQ0Z6fGxSED6+VDV+SOPC6dhvhlWzEAoOJkX/V5nYnEKfZugdyshTFkGhbk/QkRKMc2WipQ3h30y
VTiao9QhoLdXf2jZiD/MxCqOX7pbsZ8x5U6SMYJBvv6N1bL3fajZ1LIZvpsr9abwl6Lzkg3XPAEi
H6Q0a1E9PZGqeAEy+ZWktYFO3iieZScH271z4FlDkreZSqDNnJSJ+G0eSKf/8KsS8fZITbRaLNPR
Sd0wkkFs4AHwRQI7sLauZdNvu1yV/5lIugmPVyHWGV3E7ga6mxVf3lrCVPPtoJ8JZ7kBy4R3KTMh
pZzFwT5QXcfOnJxBlh/bK1PC9zhDnbPqiltmke6WXIsFXJCEThxKy5CP3t0J5dyblxt26PPQwkJX
RnTn+nh+u0VJRvRV6YwaPr7VKfgT56jpHiRg5wjand2ZXit8oHgh/IynxsLtrzdp+KG5pWvvl4is
R/HO5MRLJ7w6H+oukAi458k16dZCS/BGwUmnTNdYO35ySPMs6pGwvLKxkZHg2lINWblK3LUHcq+y
sL5+tu9X2KXwiu4MjJM1vN1B+N7YjCG3j98BeApwMWsXFZQubFqMf7mwXw0KyAiaekdKIzSTZ7xr
hsOI1758UK7bk1eCiIBA1m2Jp2Td42Wor8fOaOkAnqCzXyFNZexf2wKcngNrI/TWw9U00VCO7bHI
tekxw/6u7WJ/alDKDk/bWE+MUIPe0H4p41nu1ZQwyJrN3qlwfsHYQL/lA82GTrTQpqsEVnqHyTAy
WtVI7gjFJ4nFpq2xfGPtOP/YVuH9GoAgYOmIubd3adfm88ikDXTEyu0ENahVWr/VRllRERXDugAm
R1PpywAKTw94ifvUu5SzSJGQq3yw2Tttkp2pYB3jNIF7IA1jQP8hZwnmze62oJwDadoxdmSs9ul4
YKUUqRFyWZRQ7q/48QL920maGpxiBzEG+oyyV/WvH68L18p285nb9nXk24J/vOvNmB9kYFdx4lzY
3wfhOFx+s+3WvLjggXZw5ioMRnRtdyfCb06LZG8IPn7135Lpo6CklwLOC2cbdG/BW96pPhIWy4Nc
xPXPZOgTkp7S1dU7DZhuGmvnoF38QhdwHzau+cru34SMuhiKVni4WbsOtFMdgmLYDoY7wcDzX75Z
O7R4tVqNq3CXdltnYefSSvCQFJ8Rj9bRgHqWPy81SbTVtWzVKZ6Kvli23Y1M8Il8lt4ynP+Hxgdj
xIIawXRZx4m9cnObsVNA6a3B4NK00sudc9vs936VBsgJMorqnzzB/XkgnBB6KUaH5kgC/EyhYyJT
DMsnS8syTkTIZhk/X/vhXNR5+04gnXnFkW/bWBSXhwv61nOYNYaH9SSmJT+eOZ51SSgWWQ4RQkNZ
+t0WjBSuH7V80pOR284NX1L8Vf9lBuJKsnRl9ffx1oTlzVld7ef5U0+YO3GwSG7urWHrYWVeHQoG
E60nJmlUtShu1rackonk2t7My2cK2ti3XLqzBkFUNTM4kO3al668TwxKMzt/zo3RpdODYOrXqwHE
XoYIzaxMJl+lTYNy5wfIdtDmmaDKjpyUQZQETZGMGZqS1sZyjxRoAH7zzYMqTC4JFkApIfUrXPiW
7t1b/pKp9cBFSzoOpA2CCjmjF0zNzmEHbjvKocIByTK4YFpraZbx3Oo2NHQ/wdFI2q77L3UK+ohx
ljeL8aa0R313MBTmrGDrTh5GAQ5PerUobKtXTyuwjvWiejE6gymW/U1OXU87LJM7al86qoHYRiS+
PaMtnpfEla6580gWDe0HisIZTCwxaRgan1fFpw/+xVy1EwK9HT/0FoabNi2oCZk3QePLV/BMru/J
1QvGT/CLMzzERiY3LwHNy3hjwR8YLPcR01o8KdtYeBwd4P5RL3yv27vxKI+IyNLsUidChgPFZuxa
sOPdH6lUWMvxPNRt1eQFc7T3Hlu7p439lhkjxij/ljKUKyNTeU6nbgptCzbymMTWXtHHhtKPN27W
/Sy1fUCfKo5K/jgC+Aomj7IsadKBUP79EF9oexIlSLU/Pkf0KbzMdIn9omnTgKjv0TkOYCW78CiE
fgvRbuuSLU/DdDbdH+y/4IN1KiGu8ZZ8nb9LVBeRNSoqCccAQ8++NdB9AO94wC/Y/Xi1UrJDci7z
3F6jMGenwi+vIk7iuIxG8d7QRYojCcbJi3t8ydgYYla/Wxyqabs/36OWyHECTcbv0olwjhPwkeKE
sKDOPcYwjrTWBXo85Pwm1E+ph+x1r9J1HwZNDyXQH7c0M5i+AndD4Bq0TZ7nnnSVmTeiLs1iL8/H
JCTgFJRuvqYvnLLo7KYsHPITFRCggGWeY8J1zFzfpU48HX4EI03WbEYFabcx5B3Hudbg15O2eHyy
1OuAIKZfIOIB9S3YVGebWaGaxdzLCg/MfSYvIMc4Wdyu/Be8b6rNoE4qqL/xqfgcp7kjGeG9Et/l
DgRuBEDMAzrJVwibQOR/WIbMlqIm4vzS3uLYv29ULcsDD4pGPN5lyRW6dWaynb+54Y4Y6Uh8ovq4
ADQoQ2++oQSKzI2VxQHSdD2Kksyqc8LdwLihDuo54jjh+H3B/gjae5QuIiJFBz39OuGfsNVvl43X
viQ+yeeTjcetPfW12a2PDtSS3dXGG1AFvQRQOkU6Ywb7UrJF2SNxzgoqUfoVAF74nNcbEO1LxgCY
lCeeD+78FWofFViPgw+zyrdvSE1xunoKt6HzRCgCpIN/BM0Ns4Ci71lypiIQ1dbG2KzCCkNBrSjn
pFqaiND4EMaAQGmojp7vwLv4LbB0Rd92CHEQZFoA5PIbvo+dBWTdBgdpeKiLjJn0KO/lV1FFJspU
aBS+ttmBUTHk619RN7s62DJYVTJlgd9Dxfm58EFyZlG+tB0kD02oGza2mJEISishqiHzDlVFMK97
iouq/UG6sZpilmABLMyxEaxkKwJEfLCH31CsGDSQPIpSwzpZpJVSLmsMgdNc7Tn2R35pGoatYjmW
9ZP/bIRMxHH9QfwN2Fb3mCFvdKXyIq6SIhqQjBsqBlCOvFB8M432NFs5S1FH8Cxwn/GKhYEAKLzs
aFhp9s8K2IWex3MCKz5kFve6jQ/MCSDFO6+WKr6HG9RZESVB4AEGmtkVs/uTtcUTawcq+ltvudbG
b6tmk4D7d7lJoV5fYwtbd9AykDW+iSTzOQqSqCAKcNIQOsMUgsT8tn9kjFqYCYAsmag9oKKG+Qxm
FYv9kLwg6CauqXkIqPfAkcAOLIlRj7gTUSCAy9vlPa+PrSqVta0X/C2bcZHCP9HN5fq9iHzEKfhv
wyXYV7E5Ev4OhA0DlTYe8PASsrxTAbujddg5sRmkCZoFX4bU5fk/3sz75nyRKUlDkOorzkqHpU4i
MpIvP2EO9hJTfStmdGkFbITxu2QalYu1ixJ4JSBcdduzAeS+hM+9grnyC+vkD+SF2u7T3ZcDIAj+
1gTFl+mR37rKCCpL7SHF7SR6k6owkeSt6sPgeyNFy72RoVrrzv/yMqvRxOtPLzOxDP3jH/sgVexX
qywR4UdYBMoirveR5ZB4cCqchoAVy9RS/8h/WVGhT0FcWsxO6U8Y79xVY3qDcKzk5s6Aev3BjkFI
6uQBm2Txjq0w03KWEXb/OZ2aWOxu0rbZGfISTDlK/oRLZw8Q7nOuFLqPJ+s8ZzhM9vh/7wPzqVfR
CvUtSOD1LwKi0A+QQDPEe8rEP104bplVfXn18YoPaCzVOANHXr9CIeixHbXe4pnDjP1xhJ5UT8JD
/ZkxEvQvP9mwoRE0//USFILBhstWlOT314KMGPvYBgrgjTrttOTClNstbyChU9FbXAAee4CS24+D
IEVhdmVvcTj7612n0wCvLnYWK77lvzAHiyRupDGkHg9glA94WLjCByRRorXZGTI1KyO2eIc4TgFE
ofrP80qZyfA8+z0W32EA5x16GLcI2wNaRIHZohhJiT/xg19RPUZYad0GlaXt+FElh4W++esca3ys
VIqlSfsEcwjTQd1vEzeNwTnYCK1xe3BtshekUAGecr+OP5+3+K3TGa1BK86XRktRB2RfMKe4qQ5q
FkTYzLT6Wbkof9wjhOnjYlRTfXGJOgRlf4DKa4bl4p0GXnTdi3QA4YZjF82f8Mi1OfI51qxIKoco
2VvJ9IEtk2vvLotCZRkyHC67sTjA70NbA3/9jSECK6yDkqEDbCVgLDgA7wbDG8G0RXa9Y1Bwlixu
aYB+Ymy9JPYvxVWzW3C4tDOnym1k/bheV395c3gfnURRO4CWdefBffsSZmFskenhQS+Z32p8sl1t
WRCC3nwjWTtHDDzcjjCgfBnzX1BfESTtt/sTgVeF5L66IMM5O4y111edd6PBHfZiXfR6SzwltOg5
DRJmqoCdKwWcDS3INGo59/XxdhbqGpr+5RmVjil8ntxGRntp0qNGKpWZcgrJuIiLnQ70vQ9+9zDa
qjaVlTNFViFo7k8wlcfUpcu7zVGlWDL5V0nujt8feiQwal5LNM6PWdvDMjiIVdCl77r/nwrLZ601
R6bs9j0E+QMccUkO7/vaYHGkuWP2YphoWJvzSVXyxjssD9w8r0f5wG1ZksYimCTvE3LHAW6riWJk
jtWWwjuzH0IgM9HUgWmzfot7VGRw/ZEzqhAa2yspE+OE+jIsDhkzTp4uGWLNXPKLZqNJ5/QLG8uo
y9+NJ912CknuSFyeG0IVHqcXwy4FJZTbPgqLZYWdd8K2nBC/5kQ5oZ5PJ94i1EIzrAZHIuCZl0Qg
FanLMjSHxt3Nvqp+0M1jbhQ7ZpUpL+WUHRsu3OnkxI4BPRNN/vj36NdYYu3SKgwRnn5gGSD1akyc
hEIDIhdQNZ1tIzSpWb3uEf4PKFtixtign2xgAe91tHL/tLqjZQ4qYdUbkn4CYuBYwWzBjssM2tIi
pOGoKi92NSePh67qlyxqi3B0LlsRdut47blr3ZLs9pw8g6636gTX2XHm2wd5FAvjooFIZ3iaijHX
XLZXHeoiBKZe7FKOgQ2if7k1O7GPpBioQWPNaHJOgZhkdZyocuOaeacdVuZeEA+gaYXuk/vu4//f
Q15123fPgn4w8QuJqN1FEtzRmgDPkBjbLc+/+NQmnHKFCw3lMjjR3B2xNZm6rL6tl2Q/RX7a6b3V
rxtuwc3au1WMzx7JVAQKOaoG0CXm69f35ybuzzhm2fYrjXZYZ42ZkZTVuANNULx/Xxm/uYLWnvrS
3YqVJovaNtn+rF2knspczv9VpjOT+sUdHgaTR3xPkatat1K+MEntpay7haa3hdkp/YrpIDTwl+ZR
HehdXpo9Vp0kDAESB+aDJdbXnuDieItEhfqxAgHClnBuvF27vXeEn3YvAUIVvzKp01N3JJNQR5wR
pMIR6Kiz31odoB8UWwI0HpviigGbnsSk1Zl4kLsTLBI/95As+dxhrTugC8hfWogS8WA1OcaqApIl
NJaZ8oEPEIBrLDjf42mmfu1P7hUVHxYaUCQI9+4YTIQL3OR6QxjFJHD0LZ2hU6LvuJXGcJrcYkTd
e11tKmzQBpIZ32U2wq6vNTkUtPfJRXn/2AEB0+9Na4QbrRESA5GBnOjJtK0VbMq7GEztZWdJ+U2G
5NSaIScEQXd7V5uN36TsUxE3rTdj+p0XJSYZhOIcDUs/pa3NtBhWVgrtAIb6drKJUHWL6+reQ9LG
VDYNMIMRo+fyqlAALAkDuiEe1JVSdTo4nktOQMMCmCvAhYrsLdBpoudoznzAuaKxp8dDTdbjCKjz
AbRlCPdhBRN3yGimNH833c3SAEpULUGbpxo35qoksDdaZV0Jww1qhWgg07Vbl3oa3XETkqZxcK9l
OiWzfJShpE37riEkRvwIlLbcUn++KsAkVuRNY6SJMpl6OVQr5oOf0q/sKqQZCJxRkLbr3A0Djrki
WTZ8Fd93lv8zcWBOI99+2gUYEJ8l+k6HaL/XzJayLxPJMmC3pPIRH0PNk6FVAvu9zt/ID1HgadjQ
jRBeDWIcJogRXv7lBhytj6Dysuj8BXf6Ztx2To//0YvEIR11wo6HbPozX1pxgwIWWy/h4lqZOzfp
Bd93eQeBlf8Gt5mbGNAYi1nJL8FlnnnKR6bgt8VbYsSeV3+eScMzy2ayGDtYVC0HNgnAHSVmBl7g
QtyGA5P5BMc/lb8PFfUyZ05IH4ig2w8JRjjbmaOK6mUxUxl31BxLx8X/rOVydV92n4JbbKVoZAqC
64UGCeu3Mwdy3G/esc1SjgUzqMF/n0gLAd0MddT/KRuGVL/mVCpcMXOVpZuRC35u2oChMM2kTVSA
EpJw7HrBSNULykzD1Ase6Hv1xbYzlIq/RyVefhH8JL/w3t+VmFQt5/T9+lgMP88ohDaStXFtR25y
tmerapHhFjlE2cNqD9Z/qRO0u7n1VCBfG9SBMqtq7Qcr2eXaY+iR6RjC+QgidmYLFiH9eKaJYCp/
u4nnmwbqqIiMPf+tO3H+E2XJzrGbtbM/cEGID/pN/bwRsxwRjMjxrT9CzbCkpvBElWLhUjVIQWR6
sZztY2mLUChT+BNHLqxLKB+aqo5Lpq+CoNBGRO5fZow+1K7qubDoxYO9JxB7XqCRM9M0vCBa3O2r
T646aKsGsrPuJqrBnQnTfbKwbBR9XXetJOrA/GXUoW14TtFQMteYnjovwaTvEqmnWi07c8F+p2xn
nUv4H3epA40Chlgxpu3LzLW4eD6eATa3FS/1ASKZ/79HLMcgwLaLT5PRnOSRu9gH4BSkrmH3d0Xb
mFGy+ALAlS7VIR8VEq2wxXq2OuXeuXY3DGmnvEKf1GNyn2HKQ7Ob27hPjSbcsxr60RNTApk0fLPo
WuCRJTQ0mVjBcYbAkzcBxHXppVkZTkSKsrLQj6Z2QAsVFK+cg4Aq7kXEaFGRRUbhj2JYvAGK35XG
yrUEugWAS3daeSUFSq6g5Hw8MiwfkqA1T69ja3IE5kb/WVyBcfXE5mOucbU0VdAwUGmCer/hYA7o
Dzr2ACkjfy+aVpodsypEdpnKb9H+Z46JsU9S240QQKmFkarut6iLB0HzQtzhXnnRUn/ynQFtB7YK
jwqVhZ+IqLp7z82da1rmxPbHVLIhNSXQw/FRBtaweD9t0TE2FWqAy8fvINCCJxRcSGP4gpaSBR8k
ceADV1HuArU25+u24/9rdE6qDbXB1maIkK0BJgfHvmlPn1XU6XKtoO/YWSi9H1gGurC0IU993bjo
pf/s6Yvba7P8aTGLkYubYd4vP2q+5ZwmnQNF9OclEDzmP6WKAO6ttJjWp8kKE2bW7MtGjp9zp0La
0bDlxNGtrNiQyubJvuwlumkFMC14n95EvxvsZH/n5kjvoD6L4fOZPzIGvnsK4RUHEGN5rUGeOo2S
f6nKm3aPslR3sNl4nvjUv3IXh6MXwcp/J94dmyFU9Dq0kt+QLlZdGJuAWEgOeDRSLDqmOv6aDNDQ
dhxeZRrOvcMH0SSL+c+xL4mHDUQap/Zls9yvXqpYPdPwQt8j65WFEjP1T8gKvURdItSCO+xfVglx
E/GmN3JTiSZyu9whAxR3UupbxTIvgiN3XXbHEUoBkj1YmffXpN36pXZpwCTHziuDKszmq4IbFxh3
QNVjt4WZGM+svao3bcpYVVKV1xIWNrHbohe+jI8yka2hXNRLAhW475GxMXlCJIOj2wUTuLVbMEGW
NNak/Jt2prEpeJAKbrT+9Hj4WLGV5xV+4pw/Ex3kXILrk1iwvAd58FDLVKn7Snza187i/9M7TigG
Btghk0XfA0OTqKY8PCvZeR2JFyR0TNIArOLGEpqZP85TEzXh2AYd12XQdz8/LLjy0fY+zEuqeBUc
mYaCaO3o2qo1G/k4FGmYYObfV8je0QGqqHPW4YAMwNLo7VPh3Jz9raWWecDTTrUO/oeeqKs+QD3A
PHcFhyxZZAnV9DER7ikdiIgkpvur6jrb2goyS1wTVtadqCgPOcXQeh63DAJWV65jqQEdC39NLKpM
NWhm/jIvjiOLPDTr+Yf+AiOZlxSarjFXO62OOUCADnRQBnAW+MZOXTHubZXZUhLpiwbJrJshI8dJ
wTV7TMlc4KmkBzZZMDY/5YfwbaSxNQ3RAKPp/KtDoSsLwIZ54tIRqlLVguZOdknB30aiCBHVzrEL
Tn/dFD+P/U0SIf/jXwBdro/SJAdezDA9ijoDzEy/w/XUFwJwR3rCadJxNH8vzFr5dDJQb6iFXMux
92wbuxu3g3Tn7PYXgNtN8vv5dY1NeNKps8Qk7AvGc1eQeNJVJ0G7uSpThbQbhpuY2s0vnC45r8xd
a/o4rGcalbMWW09ObiAYXs5AUVA6B2Rj9R7Hl/WIB6+4lS8NACfrl2rDOfBBhi9HGZ1q6O+m0d2Q
GTqE0vdYfJhDJwx+cTPLrIuyjfMdOaaYq7QYat0x2a6voTaNu0d5pgjCdh+j1+sPGSin31F+AwxN
8fJvQAwK7MJXGb881s71hypcjVEBcejejT2JwUyA1u48L9Ic7JB+sMT0O3mJ6HeL4KYa6mK6QmUm
Gbwb4N8PPDlWZhwdvp0zBpIWjDRCv1kIYhB/2nodWNU34vmJ/nY6ZRTnxuBxL4nhKbqxXeE68NHJ
VkQ/jhk6WXaWA4eW3QiRVZ4zo6/42TqJciMJ9x5awN7WUJKVwJYtBGJu6y/ADZ2jIzbCrdV9/6Yx
+2c6Sl9IuC4iM4yZ0WM6ZGOAIjFUigP9i2znfCuKeUnaBEhQAtPUleAvXspiCWywO1EMJwIth6CW
DeAq3OacKV/ZiWgvrb5kgQOdZWgj2v6Xq13mMmWz4M8vR/oYwPLagXwgxYTPeIQBnFqxpRJu+0cY
aJ8yA+pQtktBPB/ULQxhEQGDgtyqlXcGoWHWZuF8PJo/KYDgMojjfh4eQBICVQpn/S2XPyCH/P00
BlyTIaHyY+4bvo77xJHjD7NMq8PHX+2pc7j0foh2k+ewDRaLuTTqsUF4ToBNySMMC2Lxsa4ZSbWm
8S9+mJyt0e6wAOIi+xX3m5kZqLHcDMp6kzdKIOVTIbuYq6HEWJYoxriHcN+It12m9VDXHCcHG/JR
j/iuHTsGFTtkziJSHAeKx5jNpWVDaZkOBV9VuFgssC2J7tHsRPwgH7CbAB+iVHflC3v90bgrJ0/i
e4QtrZrJbS64o4rEs4ax99k12EoSKRldZnVlx5hNmPnAjHRMZHeEDQ45hlwjCngSc4UuNlcnvH04
AxI8YWidENZg3/MIthJA8LnkBIe/HplP7iq0XIKEr6TwxUGi7VTjUkhyGE3a6cQgPUMzPKnGYMo4
tgaKQkoRsIq7EAGHTZ+NVty++2o9KNIDejYJR3zYHwocBCijrZGe4sKU7ectjSNiptkTLd5NgER6
cxhQUZnaWoXLCDHp97a4n9YAXRoIYHTmJ/IMWmHeYoyn8lqbwM9t0WxeIMzTiiT/NiMAtt1R3i3s
GXtIFM+lxnei21X+DzkmPA9VWjsGZnHteCziGVFTTawYDoM/skprrHoWMKMCYJQx1i/+REzgiTD5
H4DHt5ipIipk7519tmxAz1SSeYcL8bFRnJSogyFUXsAre05g8+p4VnXkMaNht3juRjwZu0qJK9iW
0E/VEUL+7tj+7VxX4tTAVFji0ih9td77LreB51ratpDTQAprnRp69VBG20kr4gCPaE+BaCTBeIGk
nlQU0WymwH/tLiRy916tDday+0IaRJHLeBRpvhGS8BOeowa9vweMTFu7ho5BRECFmvscaTIQVZxO
UYqTMKpNA38oYqejVSuOO7GvAen8UzGjlES4wc6hFPaOPrbFpwpxreUZBWvdaaWTfX4ohN65Mk5c
mlebtV4iN5dkx2pPjQIOA7LwiRKNF58TesxMh3AhwF6KBmNmrk8ypdHSCKh2SVWN0IbPYwjIT8hl
IHBBp/2TgPhuTZVlE6iBS9phYP0Tnx4r35WoWaQdraOmVax5OTuozr4mkCHjKDdKfmdBnnw6vHfz
QNUHmB0I5Q3nk4Tv/8gGkrn4EJ72Lv+ghO/DNutdAwYUsUxL2BlZgHzdy8ZoTKhcqIbMDtXyi5qk
RFAmtzi+h3hN8n+HV1qtlABrFWMKQTM6G1/q0ieCLKGihnuG5YurwnFJMXVgzQblaeCVNk4WK2Wb
bdyPEyCXxsmlCdTolU8+lB9HjxwrH9Q+3w3YIxfvP36+7ZuARXFrpGECeKYeePqK9r8/Eg1BsRaV
QCtB9UU+EmFedtx6NxW99/fw17m3CLOaGkQdvrYU2ZBsamOm65iif30lrhf++MA/WMMzTqn2Lfwi
MAYlwZFdCG/MHSJ1DkzpF0ml6bKzVL06CSkZQrX/987pZtj5x+wQ7YjmiXAcVIy6Xj0JfYh9ey9l
d+LKK1w0MPAVa8a0I6AFaW1vPxo+yWFwMsnm9ovYBM2x//nMXDPU4trII48pkbAtnNqvS7y84gPS
E5bKrihh023M4QHZtcO5VYoWEZvQQlfWnoNMzu3y2Qzb9MqBG3iAHuM0vArdyBOAA/vx5sIGifre
lTlr6hi/W1GDvmDK6pofBSfUyx+hli9D5qDsFq8pXuFakF0Ai2DhXKMztCD0WFXPN6RNx5OXbbgr
wpAQYh4DIyw3AegyDQ7fihI5gMLqKCCvbzkaENNr39mFkMFNgvktvxvld25GwecCcE7KZcX3SbCB
emWJnTsgw3lXVTTeAlysEKRBm30bpCArCVypyis3x4MsNPO1GEzguAryaG+jxHm8BPFp99tCwY2G
+XCY0LF6FK4M/8b3sCvh3trFvoxxN81Xe4lX3j+7Ahe34+j9XZfy75VN2nwV+zVd0NMmLEd60yAG
uoKYs1rftRg5DxaOwzQ9oHNH///Zw369hoaB53WAZ98Il2HeJjVoLoG7z/vKjo66SEGkU3jQxWoC
MhXpVc7fqh7i8anEwIoBFpgyTgomrFLQ61Fd0udc1aynXnFLIR6lZ2MXNV56CXCmdIjEjxmOjH0Z
BxH4Jox+l0O+ghSUM7MguY0CikhCSlUGg5hgF6Y+XyrOLojOYEp6kSJ0psbVl4U8t+hIhPbrn+Ri
ZDKq2FTe0Lpi6EgUxViWckfpHFlZFlgaM2sKpSY0okXFg/RjbSU+TcHhiz3mCDQ3uY0QJvhFL+Ll
CkJ8nGNdStXrMD2k83HVvxevBnZL+1VJDQcw/sYIdT270DrOW50Tj2SCB18tx8G90TwqQ/Cddo22
YeDiBAPBdXuvYeRiJ08wPpCfKadMdCUXlrjjFa8wG2Fi4UzAcvGk4crSI2v48mO01+uF3MerNp+L
NqQGa9CtwIrFrqRlXOdSAHK6aXOC2yHwYxQyhZAc2Jev5FmGwArYy8R4noWzhWNNoTJBJ9uYBMXK
OggZZevJygYwHl/Ci/lDhQBLpXeVH8NP02DfR18urYW94xjT4JCoVRjI2+3aACd/g4ExLmipKcg2
xgdsldTeFZ6Z63g+qYnhUdgi2fQJeuPdZTFe2gVJt9E/Prr0U50PjW37bhBR7Fl9whmLfREFKxsG
9UldIuNlNfwbCTRcBOZ5SydrhqwtOpXOsVITv1/Rk7+0bA+S0+UYLQE982IQjA391aMp3UILYUID
cEsEt9Wq/LE2uFkNZUK1G0CWyVOld/woobUM8JO5LAvIBk/Wjjyl/Osq6zJrYWV3MIfxn5pISE3j
1GmSh0ctBpUu0F0wBSpAkxBMWwixh1h9USXsx1Q1+nc9uwNhdYHw/QXdsl6sIwIIamxMHYUcGB6+
iOxX9OdDmHANvVLmrw4ZNsHK6ofErgTwtap26/OSS8o14iOEK8igNTZgVi+meffkmpwt0aXICZY0
ws/2r2l74X8a/x34lSGMdqbTezNp2dJWXui1PCBmkN67fGqp9lLC1ANYocjMyQjWpGLVUbH9S2Mp
DdYQN69hpSVaNAVoWS3mYRDFYDn8cBfGOShzpKZATybSGLQl7OxAE6vwAXmcZFfMgeZn/csg/hmX
pPIQOVBplp2Lgahxe1l4AwlzY/371bNYbDKgk6FQykIIE8rS1to2D68C0j5es2nLsZXhVdw3KVe9
XFQ++P4VEz1E4o/He3aKUJdZJ0ZBukUtH0axEEe5LR853bVUZi6npk9EHK7t2586A4n4V7nh/AoJ
uX9kH5JfTkGsEbqRE8FPnD6RNX2NexfCwPeutrpcnSm2k5gFnOUOHzR6Z4v7YGAYm5uWxm/WtDvZ
HIWRCxCIdja0WGKsmEkyIUPF32lSQSDwJIEm5ydqrTgW+1tf7FBmVSG3T0ohipQw5acW3epeTeSN
OfW/LD0JGEXkDrg9DI7udNEFAv18uttMZU7V36wFD7+rIeAKYWSgWuEar3UM9MMVVpbuMD/kRF96
KEokHk1vPir5ZQs2uQZX1VVrscWtf0UnSJfkpZiUD5C8LQ8QAaduiU/1pcc02MSpO9RRqMqoVa89
bLIqDjeG8+MAYRwlwwic2SzbDoRwIhQgU5XsAzN7Q8xGEhZwPz+FFZPzvmYeLsJnIsHETkl9E/+v
kmlfm4JSIiefuvPFlnVED3VIthTr9ODqYHeB16EXxA5yH1GqcVBBjNnTcaaZc/y8d1apPIB6jC2c
IuwFtKRycX2RGjLbehshkbcCf5Hlpiv/343ElssLia7oBDB25EAbdUSALmBQ6+chumfQ94nqsW8W
M+nINFUmGRBEpbxnROwy6nT4e06Qc2Bgkh6M4K/SeEP+7gqdo41yC0vjU+wUu2zKOuC6U1ScRVOz
ET81tx+cwuvqDQbT1plekdMLkdmoiISfWOOnvvBGRjvXgi4XcQH8CN0y0xZw18KlGnPr6A6GkC9w
PMcaAcW00t3+nLrQUAa/iDUVbysDSEF81RsD6c7UI3lJh5idColHGTApP8NoSZ/+PJBOLH/SMn3k
UKUfwSmyl6h7QI94raEDB9vbVdnqzjZDnfhQMT5WMa/aTa+NBkWrRjzjTFCR8Pc1Tmtcp+ki5yrP
6/b0tTkv/x3BGXM9jgSpsJg+5fsibKirkPZtYn0mEozYXW95iTrzuGN5AU0E9vQboPag9rhVCFet
ju9gxJPKXv3lM+82oEd68/4ONyN6qFrRmg5NughOM2JfbxIICJAZdLFvaPH6v3qMafJjA3LiXKgt
JWnLdMHsR1w/Tk2LENNjI29era0co4GTIX8gCLp8gm6CbI8j+usjAiASGy1jizbW1PGBxgH4b9Tt
PrkXIT8CEzVUHjCc5AsJky79XzCqq0R0sIY0Kbw+GWxelrb7Q7bTIox9+YMadD89jF+lWzaU19SS
+6Xs7JxJ4RlM/YIGzTWYgUM9F278pJRfdNwsRazJaerlNUhiowzLqmSnQ3XRIkm2B46ETJh0ZOpk
/9fHf0xDBXyhb4f08YBQdCWUmBCf8HrNzagbtzDmnrdtKtycRXvguV+RUZJ2Do/T9cA8jrjnK2iK
C5JZEOTWrnF61QcFwLXwq57Mvp5cpMNTzOaNb/oSNZun2rjwp/8q5tEo+R6JCpR0SXir7VW2LEuK
1lHbAf/ohU7mCsSPjVXtiLlUQS9kwA0fZBQ29vGJrxypk2NwQhs8BvZh/blaNgfc6sNy+XQ5mEdG
yu0y9jleP1SivD6irl7X9qmcLABfFdnlf/GpXFZM1GqOQWs2/NG7jnVdlHKp4Bm1DGXovgQYdf/N
epVXhLg57+3oN9E6SFKwsFpg/hKA279pSQuVvg5jwCh40hMELsXcxGh3y45Qc9pVzps8nXcvHKfg
rWZohBNRXG3CYnPUJUhrKnRbHAYiRawHSJOf2c9yX5Jtm6933UlKQtOst+/mTF5jaVTyRSWFhgnw
GA1TrfsIIt4/m8y4MsvLTkBEIbEOd7QOBSZQHKlVxUOSsv0CdpBa8rYW6TRW2pKmJ685yW09XeWj
ICUevvFltVlVeXzU0ZdNb0ZQnW/sTmeaCgIJIRFevVflwyVfy7prhPE4g/COBXW4R6vMH0du9GBq
jHIt9A7w3R6/OKDswiqX1vy+HXi67Wu4LiVo8M36vW8WFsFg2BKkl3ztVcvGbhw3ZLGCLnJoE9pD
pjPOJEt34VRth8xE7z9VNwKC9nJoXmp4pu8eKXhnU2Zz9eehVXvVkXMqGjMbP74PLd/PpY8DIz8t
F+/CU7EAFECy3Dne+RmqFQQmWYnzAnz85MrO52HSWOKTK7ChSjO42QqZ6LduMaSyQyhEdQC61otp
4uDd44ci6j7y7EWykJ0GLpCMebFhpv7YfWmJ+Ke8zmjp5xIcjaEynDjKVZJITJMHAlRLjcc6+lzG
1bVuJZZDzF2+++ixcPEW1GScu047djb8NiZOL3mUCK49VNmWTeRuHeE6oI1sVlDWSewRJJlIPJYW
ILbZw0ErnI9ZGJLPpU18LFdyunY7Iuaj5deIayNNuB6bNQXVzSNMKvpK0ZwLVYFb+yd3qwZ/9aQQ
7VGHp/BZeIB6+Gut/o8tRHjOhL175XTFhfCmFmNkPBpJIc39kRJTeSNpCiv+0QthAc+DoY1Kp3wc
YdfR3/Q+He/3GrtD35r8wqjNQp9J2ESElQmLZo8kSO1hZn9f7GD9tDlAxeJsLJ9ZO55l5X1/H7Ug
mBv+BOwdXLow8+SVIVaBGUVfWPyMSV6W8+2Ma874Y0ysMJdNcG91/3ZPD7YlCnI20IPf2/aLfI7V
w5xdsLxHqADzNV6Fj1JPQiILKRDzAK7otd24tCMbWohwuZubATd937piyqsq7/Io2mhnkjs1h1+6
eV++kSFMYGD0LFFDOPPvcwagAbcj1/z9ML3CuJIO/0s3/rfOLyT7seraNqgCSClCCP++0pDtqSk7
SmONn/1aSub+9gMZZv863xHlYpT0OrRco2t0Wkcmq+ooYlnndY16u1teNHoilLBoM3p/x4i5sWDd
wfFosefa/h54ABs+tO15FP8o4qbx1y7jqJs2/Ph8roT18zKSO5J/yMYawQ3DPoFNY/E2nCfdOIOg
QgGfTA09ZeAUjpmmtT2caFmeGs4Tp4jQdgP8LR7T4nBcn01Ab8KfGIrvf2mKpJmeY82iGj1tTY+H
Rx5hOflpJInkC5M7422O+hrtbxOR0SU7+AR+3dZn2hc7/OfXwQEAP6l1qzTBEy9uGADSMZvIMiPL
xNG9DWmNdvLUhWwhAnf1krStrI3x1CZ2TbcYCLKJwRGFCQ4gKWw3l1e8VBcI0aumza10C4wUXXv+
Y745Va49ixgAZoSOPuwKoo3NHsC7IWi3IL9Ig9FJPZNCWSWElM//Arqjjld6eQ5sKvjHZbnXnSsa
Jo/j4XL0pxLBQI8sYogNTbnWpPsm5BftQkPMq8uz2gobp+zB9YYzDw2M+SF598rT9qnB9YrYYJsk
P7XapbEaokFVKr13oxJ3uBtetircQCV3nP0YUAlJinsgBrC3Uo4CXbZyhkKksNfXtodS4+Xq26ge
IL8koVLMu96Ap6eVLDe5ZHWWj7bs6mP7s2hOGobDqZqY4U01YtBoI2KcWt7mOj7tkbiPaUx6tjJe
JN1WAznwfN/xQzPT81KNdLnvPYu4yECmxubZ1G75O5ik+26CYOxKr0xIKyuhoEQpDFbQzmB1u+sw
brC9Kg8+5dAu/wuB9szWgAXJC9Xoi1vTJ+lpUbPUqwLqT5G5RpNf4OLmuZz4K4RKaa6UKeDxXt/5
SqALXGsnI5O/+4YPaydOsXDoYL0VkhEFamAKZyMP251nMtRGm0elaO9u8UPu0ICp4PC7G7xvg073
kAhnkBP9T12uow6i64YGsUWTzcKy5+IYs7gf2zzIkm9+nATo9QpYxekjt4AP54Y9DI0lbxwF03Cu
DYAfsGE5r6uhWsDfUc5NvjL3NWf3w1Et+XlWQwubypzqJqBwFH1xH6LrKI5UD3XkAJPERL+YNQsj
v6popx0DlbWO/L7R6ZfNs0A7mofaKW8dLRbKHQ4tFg+DjSQnWpXRRbCGCtHZHjtm6Mv1B5WnrbSQ
8MO27YP/f43u8z3err6jfv+1E2QBvSeq76qBs54Ba4v/2elg/OBJWxZrEA8t6IrRzBgugWXwQ5oV
x4L0uyQ8ulmONW3wfnon+wBFmubuKZTVotA9ArePfbzlqsKMmhFLvlgnlavUOiT2MSoMEoHhl0hr
6/zAscgQHdoXCIArxeGv5FNSKjXdOEr2u6WkEYh7f8PI96bh4LCwuZIFofggWOwXeubSwhoh6MqT
nzIIDDEvEaCp9KQLb4ezt+f+yfP2o1C3TlP58yLqc3nKsqrtVXwSwdCccepPunG8nYcOykNyOyL2
bzU5rVjtVBXlS6nrgt8a+LpmABQKG0R6DnT66exOL4fqv6yg3fem0njYa0KJUMH/uU5Fo3gqv24j
RbNY6aalLTv+hiof3MFr8fg2j26X+IEZ+KaQ1ty36CjcXN1/i5uv/3DKD7inHEZ6ID7j8JK7qTFV
msk6ECGtzD7kfUgmevNxJdfMWfYoEAZ0fJ58+2WT5QFVh5mpNyOhAN9y82cWhaA4a7XC2WebHvxr
6XcC71Wsske5pefuPYLQLo93g6YcLgj2PrGev0oNpcfU0dCyanMSASdCFbx4d7dC1M9wYyRdF8rZ
lJzlkd01Z1onCmHaOAix1rEt0avoX2BVPL/Q0tihHpxY7fm0UBXgxJrR+J6BzIk7dLEjHudn8AiI
NmTXyupZRWBuFL1tNQz1V7VHWDIJ2gAzB1OmUcB1y7n/HfcutVrqwuDG7BcWCMiOlsN7nxFx7Ha4
4RHyBDcvQ+GzNR04hcG75wTyU6BlHxycMcjTk+w2t/c2zzneOVqbrUoRaM86AYURtEDpY8YsGeHb
oJmSoU9FatAfr5Nuy9zh7eiSdcc1A6B9svwW5glKD5wGpSuwdqL3d7PgCdqjQ+wUY0Zopm5G3r/8
x2e/bp841cXf2QlnKAFymKRio815VH8iDDOibmSRKSSIUivAC5YDq2ThvHWf8mrIuuUrBDDGouQ+
aFVI5yz2AuebUr+bYxprwbzNfIpuLeOBWnaD/21b8XVsSWwq3ptPq2gxN7iaik0Ocf//4WgRK3PS
6EgT0yCCkRZr1h/mxinDtjlJooDeBSt9s7YlkpALiYZKlh2elwwH5uIv1Q5DiJBdivuE0rta1dfe
8U09OBNIvaJzrmLsfK8BLZQ2Zi3iUQo6Yh5RRb9iRkLELrPhbELyslEkHvKCh9iO6s2F9MgmvilN
+nRgAtRhaungzLkt+8txfPAuX7AUnIH5ufQVKU7AsO54JljdGbPNUV2W9gLmvU3BlbWuRDpduCHB
A3xCQ4VnRg4qGuiWCUgq15FpMiHA1CF5k2FEnqkymQjNhzaNiklULDxD2uYWhRdco+19I8aYbUTf
P09RRLZrVPX3bJwlYfNcQq6EN6YndIez143nxKdYIf1Xjvx8Hr/AM+oPHn83UW2WxsuYiioXhlpa
Gqj7J6yqWtv6nvZ9iWTtexQaDWjHDxIgmXNdJvrALrMXL1BrG+1WhpDZbeiWniWFWSjI3MCzilDa
HNnW4vrtqhbPUFSJxN+H4tO1DRw5ZjDyyMsWWkkb36I/Yh73s4wLWgeIbYRhSyrI3sqIBQl3qHgI
8kdYLdDysXbpfMpS0Yb9N6LxAK64CwzQ/LSX38o006JE2krSQPiJFIod+iLnsykbAQHbB5m1grxa
QQECwn+xDABqcnAXpURd2m5NmM/bDIrYzhlGDi66jVkGUfZ4tJKNH0ThikBgFlK/oLxGTnD5cUnu
UeAlxyH2qDPbUcYZdbdY6xTx764fozwlSkIs7FSOQBfaVn1nqHRvQpmoNN0DiDqPE73fWn/HWMOS
b9iruKsJGLGMKJW45DZxNxY6QRdHuFNI6GKzbVZOwHkhc9WNDrBIc3GkkGWTze2j6TUR4RLymQ2a
EIFtipnV0GeJm8wttzjTby6Ae/n35OsRc2z6ZiEM19TxxxqcuJPMi3HvGblSNK6w3/65BafZWh00
SGQQmMKps3Urwa4Bioalz+gXwG9FxL1E5/1xLdjkBqAWPoumCo9vvONamZ6mAqU6etp+VHhdcK2c
vQQ80bP9gB66b86nIri0nZDr/riz55UwJTtrmImfA00EDJa6C2z82JIQDdJ0BtV3j3QNVDGj+UV6
REfo6vIKEaPTLN9tLF/Amj2oJTfIt86cZOY2FgiHAhmRXi3Uy5CMIdEE1bI66h/tt2Na63qJxiss
IedqLBYhZuQnASCYE6fq32b3WPeJAhyFEOUQwoL91PQzVq2rnD9FQu7vo2HYFlKVBpkN2HQFc3Yv
o7sl4WPp2PRtnXrsdq2/40hkcnoCdg1Jt+zZZsgArIWdpmYrjF/0MvyHtf7fJU8qRtEMyXhbr/0o
OC5nqaSqin5eFUlQhM+bBHxqEB9iytljWUjWQ72SBaQQb0NwAB2KiHPrkPz4lKb3JKSfRlbljkJz
w4vKYyEkWlFTV72oDAdkqkAYKoAcp6V1kmYB8weeeFCTtnRFt4NTwxWrmRv5nyUAgiryHtedhzHa
TG9lwfHPxa45EMddj9fQb9KnhXP30RyMFxkqobHlL3SrDoanIwlczmKJRaY3mdyKE0SCNd20OOtq
NoaMhahwl+2WWZB1NWBqX6ep3AzkIZzhbMW5287WYMSQBH85m+1e3TBVyxGVKI5+VK2YwL9wbkWU
Qopd83zEuPT6i/6tYlHvvTjUryWUDk13rY6Z3JocvFqBkvhr+e3dyGHiZl88eK01TuMoCp8D0/3r
1dzWuJMC4HGYfS4t1ICLpejoZs/ddaKYcfjom2gzBA4eG+3aJj+GnYBM0wMf99/tl4TqqBHznPX/
I6UTECDckg9I/l6B2E+o5ELw/E/RYrCxuQI4AI6PW/wj6hr7JMeW6WhtfMmkf8bpVtR4mursuWhQ
eQtiKIxuYKscLgGGtsc3dbwLEApX+3RvSYbwSKCfq8dIuGtwxCxBel8RL5O3lY7GKOGN3OZ3S2YA
u5q1O6ve2BbVC0o73FVyTrvzmxwRnbfw6Ye8S2ja8jEB7rM014TqP990a7K71utD06lpKk4NBBM1
wmdXEgQl52KjpLGKdJ+l1cFBAJVS4y+Fh+kZu5zFZ8T0OwVFX5B2TRTCqneb3GBbQFcTZ+T0G4P1
j3plzKYokWZYHBkjjyqR7YS8V24r6t1R+SWerWMTNPUjaYC6ZDz55rQD/2bLcFXqOYRJQpXU61c/
TWeOmMh7TDvgOelN9S4K/6RJGKe1FnkUBNMJf1df/Dv0FPJw0GK7wwqKMGCr79+XnMe3IZURA8P4
4jk0W0Sb2chQoFuQDQPnccfTy588iJE4pH2tFlWlhQXYo+Mw4gN6i8CsiVjumji+bDAEIQJv4XZP
CrIFSCeq2gt5cmrdT6vVBz3e51hZZ4lc5h8aWPqUxDLm+rnZVkVeJCmYXLjtsdsIhOjds5NRyKUf
HG3a3IVcv7scag5eFCypBRRBKkxtlxUdlMD4npEnx7qFJzFo6nUb7NWkMlIBS8laaMGm+0WlrqvY
hG6aVkRiYX4xaq8oCJqodg8KaDwlR2fqSwcF2aC6uHjtDCdJmruirvU+iPEnGP7n46R4pkJ6mn29
k5wffCMpM35k+qjfOAhi/PJKSXfYajeBWqVyr9N5l3W6u9D5xzx8GejJSAoOTdwi0kajoYewGG0K
F+FJ3F7g71q4cYoiLdqRIn1hUCN5KwOi8KQj2fencHUVUg0mE9Bi+3koOYHK1/Hyy5PDxoFuikEz
AvIrDVwff70emPxbynbUZs0QY73wDy1viZyHZRmjJqMjhwACVzq5aEfktJJiRD9hy/E3l/oOAzNx
3Rm1vYRhG1M/UNzRS/c6IuQSTi96gkiX3NUZy4ESkgIUaBsMbroLA2vb90AGY7N/vHxRvKTlmEL4
njeMcJSPDvlAywTtgwqdy1BgfrrRebItsj2TNEB8sJgrp5g3HKeQdesWLuEQph14Fak2M2chGbZJ
WfwEPb7VWWWogGa86w//D+MYx/CkfnFrMpXhyp/TwZotZTLJBXZjVK6ZyA2K1rwVGwHlqHDHyS8C
JV1RpCXYcpfBjV42DMgxZjaf5EJFzPT/a83i8yumvZdetJU0ErhDBUNiD8iS64BOr4HeHcm42K1w
g9Q5KQ7Jl8IfEv99gVBFn2MUE3oKGEA4pQocKL7Bugmfb4J6M5zrUaMWzM6mzL1MpKcEOV66jECI
V+BY6UnYtJaWYM+D0qy2eHT6NAX8oCk0LQ4F2EqupLsIMiUIuC9apexU+4W6x5GnwvbYf8d7Guju
Iz8R0F1lNqnTPXU/yNPNFW51yST/RfJ+k3OfyzTzWj8M2t0tEVxABUoQSYVb26yqPflkWXB1/96l
hqEwZRQ7Fqe0qE1EvlZcCn3zGSRbMMYSBsoRyPu/oFvhVlOQVB6qAe1PXjy8hjMapNwiYQsvgsR5
iIg72ie5So5mihxyrbUOjVA7B91BW9jkd5xxoXETdS6j7qwtpi8Iql7BBNRSNjMamlAUd5eaVmA5
EWSkb2lMMp05ilmqOdV/Qw+mtJ9WRlQLhbp4cE/CmSuaMHMnQHaq308HsT5c7HdaVsg8Nzc/A59O
wiEZy813r2SmhVpAYU3trU7L6Cr81+FqDEXJYvfOJcg1aWTaUrzQwYZGPV2yJRkdvZHmtViaX0fn
TTMnt91CJK9tcLCHMGZBgnX9cGEJQtfFPgwXERu16YjdbKVwWtu0y+OclotYPgzm7SBRr5Wimc3m
MlODYlSwYL02ldi1AsfeE220DVSC0WXOptiFC9ZeKhmA9t88TO8CZMdCIm08rE/gruYZXSgBgulN
6OvoTeUDlSDRCdh2a9SWH7DabyJiDyPCJ3k9QI3g4lk2CIzQQO9dKYXublI1uMWwkXBnZV+FYy4K
PxdSnFGwWy84slChypUf28UKVK6hgcqTumL0iR5S0JmlgfM597hc3fpHUpeojlBi4APHHJNwQx/J
sBm5Av5tfgC18dB1BovgH0Drk3JDlLREZc22H4FL700IGShvxKbO+n6PvpweEPprUReB5hxZrZ6X
8OF8fnhBhYz/OxRosFOS8OLUTW/vsea/HgAYaacyAjAJ7pnKVz7+1Wnx5HGGH0UHlVATIAnJZ6yv
7U94IlmC85HB6APSSv8IQtpAH8RDm8M0IT85xdb8kn7g+vWnTDyUalTZNWfESwdwh6OpBHDwL5zN
nBd4pBJ0D8H+XEdCcV+gC5GaM2chAGxU9l0KxSIK4Rd3N7/ZPKdIKQ41Zlzw8oCE1JXxVyCNyYcD
8eJjQvTR5cbSz48MBQPc40VNe8LR2dqFOtfZptx2MkpNUhlJQhRZfzHMsMwbFrk71MxkOOa8JzTS
uEOTSqbT6enB0MDqVEOmG2OFgMxLkEKmM0CFCh+BCrdGpdSQmW/7ZfA1KiqbL/7HtFhutfmrgcZC
UY+o+4G3a2OX23Jj9DaArdnAirli5SBfQjDBK5SSiiyDUgxYKUTt4VOSLNAUNjWPgzDlEUQdBQ0n
DlZyekY1lHULXz4fkhyx78cU2lWtMFP9apCZOCJGzqERdsUWGY+rfA1cuuUsRyckmzC/E0GvFhUv
eLRKnBD2GwiEmcgfw6zOsCOCoAPmzIHZTOFKH/KzWl8IP82RDIjbKroRKK+k1ZZim4srBjSq6jCq
V/RBPpvYqhzSX9cHiXYqHmrqZlcSKgKk2RT2lhzlC78BV9yvIDNHpW/pddvSMXUljdYwXPCoLzaI
gEIw+z17z8xR4Trj0gU1hRzVX+wrwPdnKQeVzI+/rWLBB1gMxrYSmXTHHs0hFgDTcZphrMKqHWje
p/7mfCDuBDlfE249rWuPBJuHBJUGutJJV3r6i9iGbMU2ENIS2yqVmTyYS0HaHk4a5KUl+0jxVCIo
W+v18/DkmXWElLeYHY8OF/ZnXlm8SmVBNtww9+hu0q/BxfMoMU6yEY/SWMaxbc4WG639CrK/YvyZ
lCQEF9KZ/xNZQCRGj8kPxuXWCJGGi10z9QgEErs3grqNJY8R3y6wLaQ4JrcT8Pn+I6beqzyvHP0t
KAtlqTj9+p6huaOE97eZwDsSF63JrkQHS6alkTPKzUUtVLYA+VGnVVn8ZspP5yY1vM8tGTKPRYTH
PtcTSE8rCiJqIzPkiCeL1GREMyGG8z8HjbKf8qdSA2jM2Y0/qB3SNUYrs3bp3CXUCc9S5wuKbZsI
Pe26UudDURoJsKtJnGhy8TxaZghqJldBQe5NZHydWV8jUm5BI/iOWKUn5EJTG7+WkcFkTgO3/icW
TatPCbVU9XWt20E81cm8qxoYFdLfKbSijE9UFa6p6t/OAeXtQBrwnLYvnCXwS7Hq/23DioDczQ3L
FDqHCUKdVTDDpOy7grC7LR5FNx7fqDlSCHe1UPbjntc3uF0Sod/kNoLXzGbVEpGWZPxa2C9vsyb7
Z9H3wyZb78giO+8aSHBN486lvF/NRjtgpM4D0egCanr7sy6XvFVFbZN3W1RIFJZ0NcvfZIdDS8KQ
3SBJmkNQ6lW7EuB1Cm8ObKzX/Uke/PjfxlSSdYU6Xbd56IeyGV+3soqt/BwMfgqfjFNuJYbSrEBk
uu7zjXvXppD8RGnnbWND/pJ2Q9S23SxRM+hbjYey5pmkIrul9GJm2ZSO50GICHpqYBn8Rh2f2o93
A2Prayi/euzJ6DoHSNdEakC5awX1diQqQt6V8pyIwbMdMDFSB/mo5/Fp2oXbFSzWshMs0nEmRklD
O7+0uGEY1IpaGlgo4yEsqmyDn0wD0HZJu5TWyyzJPv3btc0w9xafn+FQZBIYxtBjWrTWa0ogDjg9
w1s+GK21uHCkRzCBEG0CDZZEwO6IpPl+dPH/a6b+8245Ejb6ZZ/nx60CCO1UDPmAU/HLASOKWW8I
sHT34NWCEfqeIskLLpuZY88ImhuMwkIIUbPqqyfxIgnG7WJugPvkuQUbfUkZb/1CVKrNNn0AyKK8
SDcRek+hLULl/gbQNtKtv2ehZ9ZrN3TJEb3edRXrgaN2j2uXYoA/H0eqRinoL1ZgFPYEu6g7Owme
0HOW2UDen70peRj6pf8me/lhefGbZgEzfu3FTJ7i443uqyY03JZX8RM0tI21KQBwjNVcw9ged3sY
sIlkfKAIsWO0YqIUS0QGzjIj/6ZVulBJIgDn3ahz7rhPl8DmBdQ7/TpAYshSZiu2MR7wTqsW+MqH
nMvGRuIt683ydgrJFgmbE6ZTzU8BwEFGuVeCovYqDjZ8R/y4p8Tb4xyGrT7bUiKIVYqi8tMXv9x/
sJ8Zr8FpkIuKqjqMohVdXqU03/sP22E7PZp54LEYiDNtYTVRUadl7Gki6weBNWh/Wlzwx1U+ZlMK
gE3QvVBFIc1I8rrnRIUihZRh+x2hg4pmtJEZiaCdoIBKnkQL/ZHS3OQ19dd0KruL+LHQwPH22Flb
tJwOPCFkA6oqkNMjlC4d6IXJ9Zl3VuDMIkp1887CbkwkPcNiL1rbDuWU+4p7mEf8trsicg8zZVLR
HFm2LvD3rs4fTsdWXg3Ng/kdddX0kExwUb75bWGC1c+5X4umtjMwA8U1l9oeaHejRVTrrJDaowIl
fiI0iacgRkmi/3X/k4ezUW6e0dYKbYDyvK4k483AxHi8zg4VulQNGN+n0LAM9rMyTJ03sqrUW4F6
pocDFNLZGM7D2VtX0WfTy4UhuF4AYHGjvft+kNDZ6RruoZXqd8QkvvfH5bort7nD7CScVBpg0SzB
wms1CEB8A764/2PETYq7fViR41/2ra4Gk1iF9JHQk5weDIlvjUmldfKOVXf+t4mJ2sHkmuNHSfgk
TzZHW8nNohHXrV1JlJv6h6/uSOfcpJ9Mei+cxAGGzJXQLJHcvXrudLDzVEWN4EShH9Y6SRwwAzCL
bpISCAVb5y2762AGkWFP13GWZwxGOq8ya4adcAdHEZrf7pEPQrZohcN0wsfVkq5t11gFcD22EvSA
a/i7lkemcouD9W8smKSe/tF3vlshQ9Mcpk6zKKANT+rYhhm5XJNhAsfw6n8XQgQGLd8d9zP023e8
wRVgWQl/D75Hx0TOfuMQWizLVa80sJ4NUwjxz7dYNHlF3YUhZ3+EBOulvC7zBghxD5DquPP+O93n
HP6fsZhXS5bd8l26qcF7vsyZpCmjrOErs30ZUQUGOlEyu5dAuTthKXbqcf8G9lcbr44noom2MD0g
hkYb2+T8KUxbyqAsup9knV2m1f/2nwFtJSaL6Mv5ZVOBvJ2OSyutZ5aKq09Vp4aP92mRpt2WxBsk
b6Mdv1apDAfS892LhMHiPQrQauz+jX3DDAn1kU0fD8WTsIzSw9iPtuS9ISp2xXm+KagG/8SActuQ
UnIF3OscQTCNPRkpQgyG6kfGyU7btCZrucE2b+EJGukvpwYXypip8RK+r0eY+qkNn0OrBPf84zVv
2wHLulJDgxIw+Hif2nIWsKNBdGfjGX9wlUxSend+jXWCoHkPDoxlypClFb+xKFEh6dawcTexsIpD
237P9O3ifNR7HTYAhMEDDwQTR/u6oj5mE9911fTHXLIbQVAmfoQxxXvS4+qBURrjrJBm9YdbsCZd
AgjmWA3jUS6D9EJ2Yu7cJB5nD0mDzkmP+OW1E1sbCw9Ir2tlaqy2D7pfTf5n3ZzYpDjD+vdbcpdv
TP3w7TyqVnRWSUy6Jp5EVHXM9k8teMeQfHdVM+71mr3t26wCf9wjmkQMRI3AvDj66DjDxlcy8x+k
rZ17A28OR41zSNCmGERAN4NqNM0EoIfXAPDYNYnezPcphmIrXvW/hX+uxokyL36Ci5bWbZ7Lmt/J
CcRX8eW/h54H5BnD0G3cevbfJTVTHgCZa6x9Z7OobwzvbFlenSH5aWsqfRFCHTo5vuEjwV0F2KJC
NaJiMX7VdbHnEJZRoMf/xBLbORP7VnDbnG6NSQUUxb/KYxJtgimp3e2dOCR3u2+hXpdDEFiMA3qB
kou1Uya4EP497PdfA48Y1tXaJNj5x/wDMk5zWeF9RkSNgZP2tYUw5KQjMXTVW8I52vySiKyROEj3
gKfDA7EBPBy2LiJ4ukdT5J1S+jUvfdZVcNHajvuUGrYK9rgvVvYpjO+Oe+WuRyLXzGl7d9PdPcL8
GiIiGqQHawWnvTbFwfeiBpCnscJYc4kfTcmrSkb8R60zPRw7rl/ZHzb5Pc0O1h+6wpg++18xYicG
d2GiRu8JovVNFQx/2XXex5fmHdk/5n6aoi7UUBQquNFsSki1j+ZOZ1oMLRDlma8Wqb8ouj6KoTNR
xp2N0gtX2YR9WyxFZsIigErx8PMTrTfVYQEreRwO+EEOF5QvqRC9LMWbHYSR24u/AQuIj6X6eJyx
TmoArkDylvDz6yhaZZ4gEoqtckWf8mS00KQOb1KXNQL5x4qiAX321+f/H6WzI+TQ6wUFOUyMAQw/
DLE6aMTrSgRaMz8YQRyEP4DSdXXl89BaBtbpwkLls+6thvzPdKk/2fa8YP+X/unbh3PMVfbN7MWA
pfHEl7FbVYVwqM5uK5L10pnpApjyZXP99N/M3lYyyf9+bxr5HCw4g8A8++19KLGduT9f5DgW2PdP
xBAIFdUBoCFWjD1bnwAWM2tdCRq4izyp843rX0P+3iFv4fIVeJHyTMOuciSwL3LmNVTD7JkHiIts
nZcZf9R69apxZzhGgWBEo9ioRyrKlys/OUmA8v/cdbWfOb5wc6kOwEXz9WCbrtgt/lvoRqAhjuUH
hMuRDuT0Wrbk9C1cnnrxszGn6Mhhd2pT1Q2Y/BMUexzfiiDQVXe/WFNY3ysmfJ1DogkwToANzTXG
C8vFPyflENpu29WLhcf2BnoWZiAQxVhExXrCn4saEx/wgpx/K7LXjwEdwq115eFDjvgXdvVMx4/3
Kg6G5tRtqkHmjV14w49KuvfS9fPRYsIFbJN8LQAfPOxKtX5b3rQ/Etelu4q4XQ8FqzwbgbHeTPPG
YLn1H74RjFOX6pRS3XY5sYyr0niiNZivejaaFkY/kiEmpZobIq8ANOm25Jjd/wRHY5oUiToYOhHp
0pte/E5oGjZNw+cSLwWVWgW4pO7cBWXKNwZroAMduGg3qldGArNARo98wTH0SFKucfHs07t49Gul
gMkNkqKhn62tIVudLjf7paRy4HbnWXTVmoSHkeMAWOtGM2x3DQb45Ny9e4E0Kw9GgSqGucwhKKzl
w1QZJdBURwP54gpAKlXJyvRFfKHdqOIQxm0S9k/dPy7s1PDBoiGRY7TLxn+JJqnXJl4jnfH5ZRqB
1NgjtHUMb9Vep28dxdjxE4TCMTLxYaFRMz0niG210aAwGBdvT8XNI5v+0b4zA0M8xDgnyYaezs20
PpEMGpskuCr1phnaSXEU9Lu7sjxMxJxm+JROj9hyWVXaZ+jg9+qZY32isIv/sGcgZD5wPoS3i60u
lww4MDjpDghasEyaFMq1zpY3sOLrCr01c9WVim3cayrBYRbd54i0FCkbo5Kf4g0tq0zNqiNq3WD6
ukl80HjlSbQbUNdkF+656mJ/bPEeYbD3CqX2CrYY4ECgH+XvjRyDdXxeS5qDVyRBmyLYhxKlhKYt
8TpQXcplnUxarB2lyV9VqwkauZ8nXkOacxtX1sjfZzHtYBzptd+JIJmlCQfERQ0sn2jdObS8iu1V
p9fvLZSIPd01t0BDfOoqJRGNV8Gpf1NDMvIrtVKKHN3byfoqfJLnFfN1aywQmbKvPEMmG81pd/IT
040i14UdScVJnOWndhj24wlYjNOCIDCIy/SiTVItJXn6GOxyHO3CYpUKMPef7rP6CQ7e0UWqG80E
cvIzOIx4NmCRn3HcQZtFJtPY+fxKPbq60VN5Jhr4EnOR2F7QTCu9Vmef2jioBcXYJko8OTKfalL0
8iGhhwDrD+ugXlnXf9sFBUzZPFbj5OsnCFTX7592wEylfR0wU/JvqgRV5PA+PBbPxK6f1jlp6DQl
ImVKzSpgDOCqNEn8oVd/Yifvnh8wno3w1PULUBuO1WtDUg0MculmREa6TUUxuxJwH5dpDmsCaeYL
pVrRrxwNLp9qN7G1b/LRCcjO40vDwEeNJxO5kxhzoXgpmMzgd7ESgLOmEucU1aanyE8VA/7a4Akt
hdSY3adEhQ0MC6cL7ajDud5slPW0ZMNEgA4+tlTZYwk8LOD1OUuYlK4hd1svSgB6Mqbl39P6VW5u
uw76mJYO9C4ig45Jh6sx+VCxvvcAi3AtcoJWxJMCDg8C+xc95SN5hs3E+tg3LxOYoxhsbfbdrsAP
mc7EmErq4+uUni4o4ClyFNxjnSlYihVtPQ5XXSgo1HRhs2Q0gMspqSIjaRSGHK2tttBTtG1Spa4o
Mflyj8n5ChOTg0cQ29dsPBgoZ9EU40ECgCg08J54Z5XMG6RuFTPyjP7eTouDSKdZmOr39i1HOMEw
fPBrBlaZrrz1TwI3mwYXdNQ9Zm9ze/N+7vQ1uMe/ORZ8sbyECMSIjg2aDjpWCwKJFu4DPdpkgx1w
RGC2odldK7PDs0pLzjHqKsGiY2wMPwGhEt07v1LLM2ILRKKvuxepZEPq0dS8mSVKSgSEY7UJNrP/
HLQtiOwvriT/M94hPnW9H4M0BHyLnAqMFClFd2Z0C6J0w8jktIGPWECI/DK/aZEa8G2QhALquas+
7hmmPTkWacjoi2GI+CMdDrkQ/cHQlU9OGX9/hpBhqhCHCP8jRB0BVLwvGunc2uqXDJarIShizr2L
xEqaNOQcrarKVdSPM3oA31tjPdLW1DbOgdHD6JoTeg5ftKLWqcOWnXOtxgYF9aURzhkGVJM8pa0V
KYj235XXoEhEv/I5iZgTrWadGq8/9HvYL0gCFP6rYqQkYsluUMEITS8caIVnf5b6gEQWqtW9Tg8x
nXQnw1jM7J/UKkzZzGLvLEpvdW2fH62Xpb54fItsFAW/xVKqLTN4G4t0uZKVuDpAZif02NSe4L+U
dLrFhKV0UAQe/tEZ59MTZTC3/URwMMeZizPU42eeiUKpOakdCfb+qW6zv7JVaCdWA7lUICahzTad
zp1JBNlDWxffSe9Doe6zI3x3+iq6yqfqflH7QnVQrwt6MS9dfE1hIoNYNQSovjOYjnLGGJna04/Z
Amayv1K1H7TbpC+YoX2VUAwIGShJAgkR4AHkFZUI6prZJX7DmCscAGpRDIsSRffvnLNTev2uY+WK
pj1cDQOJO57mxXZ/32PHVZW39RibeYwTtNqXQiJrTYq/uUaRehxvFJ4ocz03viM7+5h7UgdMIOQG
quVlC621uct+piznVSSMobKBtZmM1yCaLCoItn4Bo3hqvt6u45Rv+XxmKA61GcDdWDsLoRIXdXc5
oyblqOVhTSCJTMntCQ5mrK2wRh6SxqfmxoYOvwgIHBS/V7S24bEJIMZnSvt90v6KLaINPmG2tb49
4fK91Wq1nWnjx8Ie/trVc4APM+9q6y83xOEHS7JAHRO5GZHEJWNcmdpsPw/MPPANSGIk8e369llP
Zdh8Msz+AYCYE5cX90pdjKemcV1Q0IG2ApnhcJ9rxI0ECMe5mNYBdbY1EIrvO1tAvuZmq4x8KJ4H
Mb/DKtaM6D2Yty7mHoKX4LsBYEczbvhnPLLWcVKkgjX+9z5SVFYq3uWMiNd9dlb7N/IZ3vJ8VTyR
J8dDBKLdpsuMNx1JAY+urB558tGKWmpS4lXUcpz1SRMkxACciE7MvM1EYntvJqLzG0h7B1P4AClD
5QXK+ZOWl2HzHxlM5gpJvm6wtr8mEeHl8lH+lGzX1loyM2giLGxTB0N2Djc9yIjaujsOfXsGbo+q
DlMtHWliqte8BLLd3+vP8ibjMnB4m2hIX0Xdh12IwhhHB6hz/13z2vGP1g7NbLIZyvpU9D1O3aA9
SYdrzhcRjlrgQ7Cg6DibKqqmUJT+vIV/XxaL9fhh5oHCBXdmd0GG8XCa+uJRsVLwCdKli64C0slp
j6jK5iX1PYq5wHKqHoJoL5xDfwA5En1kmOh4ebjlsTdKlXU3J+nyjcWI52peiV3J60wLoPtOQ25V
kiqCuOjNI/UeBRILLyG9wH2WT9Kg73EhZG86wDJWk9m5F6J/Ro0XgTK6+3S+R9SJQYAJtG5L8QbC
7DHdanJ7180xDwKCLTec4g/kKvYCYBz5T01WIXTZqAbKljcTMMyl7coqV36elvsS+yxHranSQb1b
WDdXItrGIRh76jiLB55PH3SW3wlnEJdBKKI1+DjQyBPtM/YP8RYpmGFYvjaw9yfkgmSjX896G12B
mKTu6Ih6cXchH1pdKmSuwcX5iveIQLuyAMQ/YKe8lR9Va6PfWGlQpCECygPmZ0bGXJQuMtusfRNJ
GV+82ShlB1YWX4/tTlZ3FwQtqfm8kJs2nG46i7R4vSqBzGHWZ481MbbnCinqcfGvRiPZysAFYCsX
GANr8Q1JwDke3XzSgSI5b+GHIYMOlZUZZMpWTZGIDD71tjl1MYeWhWrWtisFVEhoEWfjzKEuK7/4
0N/TlTozI+3Dcf9A6wuyFMCLuQ9xa5XkomVj0UzddVrJ31i8LIyZLa0N0kCNeQ4vjDxcXXvfWDzJ
mB6rqVUseVBGbSK0ZCL127wuIMWR4A+1N1jg4oILY6VRpoAP4sN2icLzBEE6iC9HH8r+8x5ryOr5
v+/4Mm7ibjl6uNRfZTYSMbc74m0ooDXal9UgbwuvHXOfZjBAuWsx0a+Xnwjo1DXt9xhaKI2yMKpm
nZ22z0HqA62R3Np+sTaaW1IaN3RX8gaabVCDMnD5w9mbYMfqHQqUHP82/cp0KNGV+cYAYbVbUXe0
gLLV5B7Lh97zXtvb2oVeZZ58wROom/GzxF5sJbbaCn5N3WUPEce66IMGdYhuvUFWgTGnZKB5OwZM
8pGNXSl4iMv7NuNHEj7DMv/UJ1YfMg7Hver3TuxpltIuyydSCyD/XLv6dfC3khBA9m+wFX508/Up
rw73ZjwSHujktVxgxlo4mCKMU8ztBXK+R64EvENx7aN1NzMWk2TUhHn0mwoh44U/tS0QaGD940EH
G7EKOYEup5GmLN1eCi4Ozkz3Te7Fv9VT0fF3zDVqLaDx0O/nB8a9ddgaKJ4zWsfR6W19ELF7iwYJ
Ei5kI414XVDguILvDMfpSTCwQaCW28ptuALOMl4lo90vhBY+WQNHC+xfb4/YEeoG2nIzOJ/Gg3gw
EHs61SSN/ejkzCTXVODUk/mggtVstXvO0v0bZc05Zh4Z1kr6ZRM9k8KJOJubCjApi4zjclvmmTNQ
TfuRmP75kr8JsOUaV+TQHSp6UGhLmIQ2dmK92u5boG9Xx/DM+xCikSi25bMGnN5vj6hZW0iI7UPi
tvOuyGBmdVRPxHAaw1ehhBRGM91jgHw3d6yInov0mxs26KFckoFlWIB2aFkJ3OPUwN+/kvzPv+a6
Zm3jvVM1tSzVqxhogZnIkkZkTXeNAW5eY+xtx610Fgh7A8o83rNSkXekL0REExDt1uWYPE2GYevL
fEqYHwOYrmj3+2HVjnTP9f2Iar8QxKTHYHZSRKlxwP046Nj+s+07NGTKMVWjQnFdgDY15H965ULD
DLAHADwwgItebzXEK0bqfBSgHq0PjOnuhm0+TT8kMJe8rQ6llLJminbppTM7NoarTPCIiykKyvXK
V0azAWuSlTmd8z7B1pUn4yvMn7fnig8B/w2yOvGj+MgdQ6sk5xe6Aqi3xdEdL923z5+cH6bHeblr
KbY60DdOzuRg7P3GWNPninIaI5UouIKjTspzO4Y+zkbBwRq8lZOinz9QZpqJt+oZwWEzxaSriCtP
4PQ2CQIgImOKyMOuQj9bRJmrRp0HmtZmvukVg4/UhVhPmA9P7w3L9mEYvUOK+7zDRQCnznHlC1Cz
r5vx6QExD7HM3mBcN99EenpAOwmQDfFXIZyEiNl5KspafWcAIKiZVQJHzkOsiH2rdLQDV4Jgz6q8
ZaJyON6gKIzm7QyJu/JnKus1vqLT69CMhuR15GPcozbUYgL5jL2R4ScMJkwEsJi8STmQnLQMKhHp
WttIspFi8qQ7pC2T1Mr6G4qy4wDszVLRMrsUY/A7BmxDKeYZhx2s+kEnsAZ3eHafbVVaEzxj+3cc
TvC9wkoyrIkbSzxWhgsBQAXwqRfN3NcR5HSLwXAihlnNh0H6YifhAjVpspZmXTCjgz8rwQwh0hI7
F5jE1lu/a/xvM7iSvqmXGDO1oZ0c9/RUGP52Sy+hj1kPAq1nGiAwNxe1MgGeV2/7RiIOABHmhvC7
A9JoeFTAP3DEr1mBf8cnl1N2EVECXEOp60cJFGDSbDRG5Dwqny1uo6yHzm9+1RCcb94bqTPrfp7S
lkukbJyV0EioEwD7kOxqg1TvNggiTwuI3212lmRKbZ4deZ97kTYS6YvQbeWsFVjSono1EmMVkUxr
Caa8nEw4TxD4/B0b9zzW54Qt1w9DiO9k3SN/cpH2kL/wxniIke/Hw0YdnRrdtYBD/tSXBbaZ1rwZ
uEdoa/QLK3JjUZkCrmussOjlCJEb+sLLuJdEQvYlJkUvZcGTbiOfW8083k0D0NvtZyagJkLzms2B
7uL61RohY+EPaMGnWOKb6YzRrKkylx0f0Mvg/JoY26+ZK60+Vp0bdcQGmWcnMHE0ydvg8HPa3Nef
ouNA9iCKPs8zp50LAepbVtxcB1AB6DBjZVIbPEtrv/VYO1e8nq0XykbkbV3BHRzgFoCHNDHG2CzS
3ESXhvVf+tUCRtmODD2fz57uHVP3m9s56wsJXmoHGtY2Hezg9E+XQWm1phoM1glQA4XR63mHo0wP
BIvXtTyEOoKxkj+9mcyWN552Ew+OlK8uQGNvviiKb5Oz8Ui5ZrWIt5y2TAYSC9k26TKBbuIuWRIi
bVSvRQkcE7IHQvk1uv8zqr4PUksyhbEQOiK8EvLiEGhVyCLyLaAaNShwZ+uDPpswWDzrqiFYkboG
XoEsesCcdWj1mXgs2bGFJmmGsu2cPtjqFPnsa388npD9IS9RrbHJcIKC/6+T3xO7MfdlKHd7HXgi
vMHH4wLCQ8ZJK7/40fIMb1WTVRWHW9BH3+rS0OxZ7lCnNL5weyrIbVdXI6qFAhbWLlAL7n+aG2ep
kESeyBus0LyjustZPJygtgkAVafHQ+RE9GBzZh9iN6SM9v+PipgIm1RELHNb9PwYmqpo3tYnXkaj
qln86GDaNNfEXARnjOy8ThvurG04fsB4eexBYvfeKo7YGqt2HGkzO9Bi8ZQg+bXtPo1tC5iinMmZ
THpx9sCG4j926RZzFZxeiHcDaGmn5YgHYNCsnjDkFSBb77Kxwee9UEF52SnqEqqKMhBU7Dv04qjy
f2LRvGnqsUKM49ywKr9dav/oFIv9lC1HtV8DydViqhMuJf3ajjBKQwwN64UJvce9r2/FYEkfdZwl
pc74+DZPFHUYrv4s2nTmSm+W4m19V+Z7xUSGZVkLhpdFbq+LaNg7Wr1iMRizR/AhHAw7GaokGrNb
ukqDGRJryHRZsEghE5bCo//aXyk1k5kGE6QdMo9UYUvEmqAgv8+NA/b2qw2CjT+oBP+DDjuo2fIi
R6r9ZDbhQaB/pXa5FScaH/RpCTQz/b/jv0Q1fkKShdK+HGXSoOw4Ub6QtXLz4EWzgAY6zwVeeLjh
f5QuA+405RPEvcCtHEq3FfK83jcnD/5jdO6FXcEs4vwQnTN8FkwNsg//fWIjQ3hWkd4/ZOLYYOq6
iNE11TrP7YM9vNHskjNgjGZ23hgqhs+O8RrEKkekeFnO7vK/RtkXr6hRw3vf9niXE0FAZbC0VAmW
gckdPtI/QYpa0TTmiXoD9PiJOKnEU0cm/JWOANvIO6QSczowYbkWL0E03v9ariXCtTb8BmEKbg5x
CdAZrAFR23lqjR4M8oeJeK4L0/qkXglrBGg5NZsJYbacLO93W+KFLQ2Ec+wB6wXcyKWzwehYNEhP
NCxRY3bj6OFg7nyh1LxDW94BJjE+GAZgCoPtPMZee23Aom26d5wxNugHt1SljjQO/UGeFfm/CO/1
ukfcrvf+QywJr9zNOSVsk5HhnEqN2Re0hBNqd8QxEYIM69Fez/ByOU9LxpLaCxA8tXMsqVx/SylH
GMbN02UOYj0AhjPWzf5NTEBCPZ/PwY75sP9tLFMyTT6dNzzTPS8sHFBIeuExqAU/XJNyzLBBwHwu
LUhvVWh+kEVW2YsbFygcEmkdZWKVHt7x602uXfqjfOzmPMsnirWm/owkn76843BYfZPWfABc0M07
7sjLE2Rs5PfxpYUGgVtwt0GQBG5CqPZ18OAIFSoXXYE40XKnSvqR82SXRmMTxcNvFpcRPENie7zl
98L9PFE5zL9rkbW+eCC1r4gWlG0AbfLIbhD+KZFFufaPFxf6BCyQUicjtrefukkapmJb3OIKQxGA
+ZjtulR/ubtmacSD3IrNkhMS3se/4bI0jWy/5qYxWlVgCBuEbtCU9W6CqKhwVEYf57oXwYOWrHs6
gZC0M8i7QQQEeSAVK1nLivQXMVVUKq6O+SbtEeDweIN7ilsKeLnU/Nk2pI0nSqRSWeN09Th/QpYl
70BRfVal8pSmyRxGFvYZcVlDXc/H8cXjLvX8aMPereTbrbNB13oHh5zX8PwXkwhgRT9tRPaG6zwD
0udZOkTGbXJ4zkQQrOc9xSOeApvCbEiX61mLL6CX+bi40ARilBdY841MilPjgfrYAqoIQiMdE8ZW
5zM2w0wucIoBswRPojBycV0er1qiuJrg+wGQGbtU2gnzpqk7kTx8eyMEJjFZ2miVFe3SlJs/JTcP
TVxNFcOf1k5AKBMfXDAuzqSGyZSwwQeGYO9/+NaESmmSXOxaUArY+Heh/tXXYB1cDdJ4OgE1C6/o
ZqY8KlDbm8Ala/XlxQTamCwnrmdEZZFuVCXCOxZLX4QnDMJwYzDOafj+VfmH4kOVDlgrPoXHT2Zj
jsLGhAFMVQx7aaQVGqIET54LcAjtynRo09M4vw246Nunw1+18G//UQyf7xwcq31smcheHOYHg9RK
5JchTUu0jNLKBIyZX/eXI4OZ/vEaDLdi8ohJKQym6VVKMJCsg+VXELORid9vFP23kdAWhtlWdrRj
kzhXBv/qa9HZf0+kUP4Xyzol6dmP0+5JIgd+cxAGPrwxdVdZYTqAAyUvuKVyUyK1O2dl1fFitu7o
wgtWNkVBL1Ou3JeFPF2N0KgbLjx9bbLV2ovIZvJMXCLknJ+acznbnmgcxhj0l+pLlk67KojauMgh
yJK4ne09RkuK8hFintl582cL1d2gWUW3LuMJSe9NAzW10wXHX/Moj2k0a6jb+Vqusqhb6/ooduYt
ykdGeUGeoAa7qa0YfRZM6OAfGAt7RvWTpMzrK3m+2xsdgpZy+xvxWwBZFjv9wM6/yDckjbArFpEV
a2ERxXUhkx/j0+Mjgn4CE8dG1ZB8WlPwwkk3+nwYOT072LsWNavPCktT3mRTaPgJFwLBtayrxMdp
0hbO/G3IEglg0J/Ys114NpisLTjMZ2MoG46rH8f/MSZ3q2nLxxsmbFttPveOfRlakmRINnyw+CMP
uTFNTITkmZsEnXyNRQuN19pMQAZnk1f6RTJjG11TASsjnsjAKgzaRsm13Yodqy8dWNZzPYsBdyRG
8+H3MJGlML9OH4xPdMq2L+xtzU2Tg+PDYY1BhxTERbfior7wzX0+7k/w802mSiCqreyUpFiQO34i
gB8m+ZxNl6Qlh0yAde4FQkIc0tCaN2rCAQMvAIJ6ki93cM/z4ijM1rmuJJz9Rteeu+3j6NEzMm+l
bn22Har9ZTsbJTZGn1H+46luiZgj2Hort088CzZgU+al7a4UJYeViZcFIamLe2LJ7OAh6GQ7TsYL
WC1pxgNqOiKqdFMFVBlvoooryTMH0qlaETqvhKNzvM4DsZNM2reiACSG58xqJovcpmatABi1rgxC
WDzd73gGewiHFpD66XJPjux/6e7rSCDTxDPNoromW1pop1K1dnoVHl97GvWvrttEujjoscCJ5sl+
Ad07zf4lsIkCdSkjf44qcLueRETTFKqL52LHTZfUsx7Oz5cN5XZ2ng9CMKN3VW8403IOud7jEvZP
etGI4YzY1Nw0++sQz0YNPLLqcXiSbGXUtGquNfdjsaAMtqHs3KCXNsN3jtCaqKg0qRQqmmyWxdbF
f+oW383EY1o8wJNvcNNKdK73/T3RPGSkGgp9uMbAKrRje3WvsCranEW9zeTjhqdAefIuORY7Pm3L
FmFjF/2KXd0TmYllH7R2NoC1Gu7jPfBW+lG10anEdHV/7dS4M4jY5Anrsn49gDZTGO+F87vZgDoU
H+bbxqunbZzDSMKJFLBHgA83ojrinbzU6lKVHk65DKhROfFtn6lmDdR3TJhYLJlFE9ea+YlKqeNu
d6AMdSjlsttwjffPBR70+pEs4NTV5+zqswpF05RExJ4hzBcICXYmdHHUZr7f/l4tv/P6UjBBLJ9r
RqPI4AOW27gyqjqxmSv8UhR7DxSVi2avmLRs8YGvi/1BkZOyA0FVS4u8e1USqtX+XyQdG/t9SBYS
f/BKeUeo2lw7pjFVWKQNd4WOA4wrekEBlfFcK0/Y8f3AfrSnC1kFjxVjD4crwni/fYrD6gmcb75+
UJRJnA4Ko/kg9dBw3HzvN7Wg6hqvewwQn4lM88fXYiWyuCHUgZcT/zkO1hVWXPK3/61gWPRVnueH
cZUF/QwRyJd7er9nFwPTfOLEHXfOwbDG5s37doRiteNQ9eesVBPx1IiEv4vkDCyI54OkeCT5bXoR
AimhfTyNGORHOw4qAcHajXYV/ctXPeQiLwuXCc0wvXToS9bL4UDSvMQ/kwhm6bhhRTw4Br8p9Sya
lNNfTXy6bQ30ynOirKnD6MHd2L2hqWBLyU6kEBBcCukejEVx5GsI4mcTaV0+NPh/0gOKGLboCtMK
LDLXj2AYgnSGOz86o4qvrXbuwmQAw4Y1WlKUtJgsZCBfUmr0Vt6aQg33Jf+fTxQEIpAuUo+4diNq
OJ6M/vvpATDcqdkX9e2fepMRes7MLkH5t2rb+kOBe+d1I7AqMBcFZg9knQapuMseK5leAlAi3X+A
k/c3T2FAYCKkhMVJ1KG31/A4unpwK2oSL90wocdreQ41uj3G4L279I8GJ3KCRlWDCroiKrk+HrVx
lbqMHp0wgRoL1J/stt+2aCJwqEhBzh3aoGI5yJleGVQ1/4AbchsOTcOyLBMgVldMd2n32MQTK8AU
qcIO+gTOT9VUB80Pk9Scc46hVDcZkbqLPE8WnzgnRvjUgqi3Ddq7sXFwbFOFT9gyJbhzb6sUF0wm
R/j0GEMNUX7i3ZurLNpIsHJBQbazPUVNH9eMFoJlv9ZVw1nfgtvZ3HYt7943XRf+7AFOZ/CZW61B
35P/kvlQJomkLBbh3EiOWiLDuPq09YXiKCmkj9UGQz7hEg89uFYvB27Tca/TtPpBzKEUtfnpqwyE
5Nn61qcLsG5PIx67jPjbk4Cg6bM6ghcUmYnm8b2jMIxwPJK+FLR4SBKa9MWDHUhCbfk/J/VClY3W
gHCs0gt0aNNTF3glwfQFgOvZUlEuneL2npWQ7iO20Rj6nt/6t26+N4hC7nnmbpqVYSmbLr5BpAh4
weiZ1bbsBkKMt9UbV54AGh34tkjvonGA9gAhrFInwbRkF8ch2qglBnOFPRZO0MjLptFxwnWjrhep
blYH2665APcPxEOnEmw7iljafUM3mhwAycEiWpzLxgwKfqCzE9iQmes/78sLHLoe+OzrxZbhlVay
7/+za/IK9V+yL7dPACcJaAxcvvA4gcqXEBIjixUnIz9Z2X479NrYb5F3Bars4DrtRNYd8fp5nZbt
Ox6oFgq6hgHpSDWrstpp8lvT5osHR6UBVLlFHqPYQEDGkcjMqWujOF+HyiyfDIm/kQJV3B9Hx7Ni
kFxpx0whj1PZ9hkwGQMC96ax8pBGRK1cD9QiJemsvi8pRuzREQSTRiAGxL0M8qS10oxjNHoFVomD
PgtAaq8CX0D/5B7R5BBrWJriz+d9hCM2UW+fHh0UIVFZiU9V77iIEHEpZiWTkMKXjserFtv/D3Vc
Dvh8c59jai6TrYtDglapiLPLYb+Yq6K6v4Bj+NcX9EtyWJ6sW3gezbYJPdQfqJiZTUtnZvm1ICp0
uWyUUndvc3e1CjvyTUPm10XAek6Dxu4+dgTMM1QM9+OB6G2e4pEh5VWzSLI+3oiieRzTGG+1n9/g
wxgFs8Zi5KzF4QI8BFIbYwNlSN6VZkU2+zefYI6hcm5T8ComO/P8m13qTXE7ai6DHBEYq3y1ta8J
g3maoS+zMY8F6peRSFCaSWfuDKWKyqEePmRMRm9cHrw8GKqhC9WfoS2pNUOSegRVjzGoKwXFbh7m
54zJQeWIb7aLf0Iurkku7/VHIyCpr91qPMgM6lZ2/eSj1beNr3qNWjPYsP+JUB+6H7FNINR2En15
zlzGlYNziKH5sPb/XuBpHj4cEqpE0OVTvdUpI7r7qaYH8MReR3RLkZnPh3ZHChRCvQDUxpvDTMzr
6qPd6ytO/Kys1c5BQrOUd0zme/kkEAHWRDRr5o/fdl0gA2ZxvWeVBBstrlem6/746D09Wxu0UAQQ
o4GyBawcjRZBdPDT0WwvDs2D1SPAvOVRb33yjbfTJNdg6qNlGh2YUmDr+M0mzDw2V3ALWPd516QC
P47vCbtbhNV1xF3Una0p4YothchWSK7wEpOPjWV+1ZF61syTu+INC68mxyG9fWOw6GfTitVoIql3
i/S8KdT/hBtO2+Wn1XrFxTBAJ+w2ZYx8fLcoNGmEPbov/bu8i3W3j7F2fqluvbYBReEc64ce+4rK
LXJMfGLdnj8/geQZ04XGk4WR/PEU+9LMmXfTY+kvYUnkzSVhbhkXCCJVtM3PHrv6WGkmGGQOAher
ddSQ30AfZwJ3KZVZoqgJbJnCjHWm0fJVesCBp3XpeAfIIerShFO4+Y/jTMNHwSPm7erWQvV9+PKr
vVosaNuDZAXZ3YR/AoKwOMD4dbskBn28PocrRfjjeF7Syq8M32PtFsmULcMgediXwRg7oIu372Y+
4iUkNUzQMYKZozxrnyBWmq9hBM0rJDB8n8Fg3tERB6ojIks8q4EE6QkXsF+G1c/M28b2L+tSDqF9
s8w8iVmW+FJlUTVQBCfSsDcyKSUfuojeA7xbT9uNkPu6dhAXqhszeEbiuiO6rHhURvt6z2WqFxRW
0bv0ICkj/aFRD0DjqTBLSrdhehiRxFM7pVCCH5KxT1Xh4qJSegBgqHIcUcOg8UdDJKSr+3HLtR8p
xaqxxIZkc9oFex7IUDKTrwamaqvmk+Z1ftfI48rnj9BIIRwnrMXdGyNUjiziDI5+KuTjnTnNBVsa
gbu65aZnWOtKfVxM+W9/Q6n2+f5TxDu8lcyXcs7dnquBZONDV9Nml43Iit53es8xoKfrIvzv0GG4
AxjVJnhalJ5udKfmaAcmXOObomSMZNLzJrEkAo+1UrMwGL4mNTEf9e1dm1JivtTZvSkxgInggvMl
0S7WJoR3aZLb6tFXBXR9xnMSTDUAkrfJiAIusTKBI3BUe63/3o/6yEmESxjMcldskcwZVhF7z4MJ
Wi/5KsbBhuI2aSpOq1fDpjEM9S9U1/c1S36d4xkEDkuTB9vjHLVqp0UsMW6RDnhGjSSvQYayRmCl
wKwDlJJ+FiquTF8ln3e+Q+R3fZc+wgmCjuiRQDHalOHroNyCuLS0qsGDORjLRwJS7hG76mAOFGVZ
1w0f/oki5NBxTtds8zOAC9Yc9gptR7uRgfXmBsUG1xiwzY7hOUa/LNw0kFOTGSu3XXGSNuebbVpb
ufYny7e9TvLxz8k0Smy1uunSk2vuTFmT3Ae+78OZ6A84C91+rKPxrm06uFZjBKCEpQdvXTFzOdn/
fh934WI5MxsbMV/QLDs1nOP5yGC3/AFXdXreli/Aw5W6fsheoe13+EnPsHBfCjmat9PRshWlp9WP
UKnS34PKOhh4uozYoFrOYUpiT9lbrylaxt4pdcVgXBA7Miz28Y3I68L5E/KMD8z8cvrOYkY6UeXP
y/NHv1jwKuZwSodDsk+hNhP3DNqe0XvcZLqw/yfFDuaz9eLIZATtxwhQND3XI7xAzc9PhOl3+rlv
G8ParH9GPJ+K46Y09xDPmDm6plfIHX8mN3pj84BpAzU36rzNqQzZuZ8/3rLQ0dnWTvFa2hpOHOjS
30Xzx+uz5dfp9l/x7QCNq0+38FYoVnXV5842nELenhz5pIuJlK06eYUd8zpz+rNLxhbnGB9zKK7O
zcQQg3FfYrayE/91rqWV5pKorlomarKDy7/igxQXkvZmIidHkhUQQl8SN89KM8CrjNYzbLEIxm5T
3bi8WbWQBDxfr4AlcZrW9dOrPC2DXMBqkasrre6dUVdbk9PwEX+dFa8V9D6riKh8dZi1kHATD3fI
Imyr0JJnBuXV49Fm4GaPJogwUUgWx5lSn0VxrjJq6mEcMyFw5AxTtpfMicDlF05wNb1Y8dwOsFVr
7MCvjvZmT0Gn0H10aekh/i7foPcKNbzXWx+ck4KN9P/69j4BFz7oYwA+3wpltVcPGFFzgumGWydg
04JIFNN9kuK0W0UdmY4n8l8GOSzCnWnoXBVIShz+J65r1B5YF+3eaquiwYHASSb6zgqKCX4JoFct
pVrISEKcYBpHhcWG2j29yC7rrMqL91RnW+rN8qrxmHDZge0U7z7XQ4hHDZHPpD8W12POQZNlkxTv
KOycV1zf04YlM4qP+vY7/91U1J3jg+44oCmk5km8f5G9XaBA67QAs5TPNO2Ck4TkY/F28sodFrG2
lDGc/5P1TWXrbSBR7dj+GXTrJMeIhijn+ZEjomyXU9jLx974iqEggsZJhnNqC0hXZYTTelFEQWWF
evEzqnr/myPmFX+3MlxlRZ1Pl8DRVr6ieD5YGA/KxmrqBmwtM4NpcvCbVUax+dgEbgyq9YH9kQrt
rsZy4T3P1BRZirMSIkI7sFgOqz/tJz69AIkbrxmFjdpNf8mFePdAQLTHJHsH2z78dluabmqc60er
wMqOTLHd7n5Gz2usqrd6Sv0/SKkOGRt+7n2CWy8N3L7WcX2nsfltbar56qTnBVZ76wvyCsF8dMuI
2aXQFVxNIvtsf3Q4KIkKbNs7hJdFfhKN3QY/amgSnvjVrtU62rX2LjDKTun353u3TqWAg1UVDG95
QsmU4WaB9fQrhGmcT9/AyEjPxi4hR4EQLEkxQ0eiiJ8AIkZjte/w8M4fJAs97ofetxHaB+RmiXlM
EyD00jEzx/nNqxq1NtN8BBtuydb3/xW9K/Y0D7sAoe075tRmKEbketYx163Fgy9+fmtR3J9L/5Fu
wc9u4RBlJjs9GEJEQrssdpYCRDyloM1nJN/dyZzm9EZBQQDwIHcbz+0r34SMV9tbLaYJzAf70poe
XZfvOZUDLGOlqUdtWfEaLjjCqvgjXRaWYTXKUbJ4SpiJPbCo5s/F/+FnOrccuFzLL30kDN4UT743
9QD5+f9XLWbQRH0AFyTHseVOyza1a+GDvcRiQUANPKbxWiKqdQkguhnhrqQn6+6UoWa3AlkJGTDr
f0pb9DtbGptOnyd3LXINP6hh39Xh5x00WWafj7FuyHZDjmrtsJKJFIFtJ+Er0Ec71XTUZxhrVzCZ
T83vp7uSfXr1cwQEI0OHrUwgGJ7OrkefQeaAJ99IVMQYJgUljQ6h1M51ONXsevkoK91FJV+ZiWW+
Ig7+2AskcCtaY6QuDZRcSjZ9R5CpoJ/P3Ze1fSYj28kyC5J8baNxBcjF3GNe4T27waBsjAAs8xsi
M3PpXJ8tGI+m3dV2aJ70/Yw/4OV9B6Ff/UdOCLFwsME8R+QR3soCdqWlsqCI29DioADVJAcLwwCk
puql5pKIvApf3val35WgPUJvttis/+Ax5Xe5CW06r8RnohA6sGbPzNPaqwLEAe0whbG+lv6b95AY
TsyssyZWsYjgo4V0rpkyuOKGVIAZh+0TmfBbDfiuf+kiMhddxmoZG+voo4LYocogH/wwd9I7wCIF
zilc5PrngiqzPRkxwBYvlCgDKoygXdDKdVVwMWYHvkPovap194c7jcp/3nqacytdGc9iG55JR6m1
Z23/HEb1yS8PjxSi6gzh6/mHAgeFOjxJ1Oc74bBK6AC0SfxIBf+gzCV6v7sSrsurdRJFVBfrk6KU
AgtpUHJDp8bdZ1Er3I4TyErnEmZcrn+W9N2JWXZwDOF6vZGDrqMqS7gGAVTLfUOPE+WCzLamTr7X
J4IOM0VI7DCz7qkwhRmo1+TqhbVpCl6NHZMN+jM3nyL1OTNTjiGB+mD8f6o3PnSkfMNc8VX+/VDx
Xsmeg/XBBKgvZL+02r6zmkwbYIX98L992kg4vnylKcfYwuXPntJopEX2LUqnkTPVDNvjoeVqoxOb
3ykDMdIv/9N9c4SJxwHakjlibbWeH+IQfGVr90n0WtAVciv0eaRDxgMJFj9ZO2P2oaNSQtEh4ZDT
is4cD+xQhCj+cfstzAybVRkz0efDICniAWlyGGJIVJ9/QUI5ek6LiVWc1OtIABL4p13OUBhQZNg+
Ys+eNgGDymfVlhb/B2NWEkvgvG1xOwHYPEUXNgDATZXytuOfY05zH/ej1oj7NHhErc95GZcQa3j2
Nk0NVdkOgjI+o+GUF+IHPfPcXhd8Z6WoN3OdBBDFLkeXiZwBRsAV8ayRn9dfmQHpSfqtm6IO0qeh
M46p14QdaP7yAhESh9ZcFzqqXh7TPqYNpjUGMcSBOZ4MTb3RqXI/HyjVdNUsO7h82aIyhx6rRVS8
bX+sX/1GLnBh25OscHrmsP1+51PmYxyWU8ENP9mM95Sw6ZxcMEnUVid2gFoFlg7BPiUvIDdS5i76
RHzkvCGalAjJOxN9yomWxwk1rZGdfHBYThmoZsnXdXcljpGiDLvhBgz0hwCxyvaG/Y2aKZb3qjqS
e7b9Pn5gbMTNFHsd3cRjM7iXqkfxTerLKLJL7I2VjdsF10cphVOvvABAJZMqcYWNqJ6o241up+KR
XdqJD+Zy/Gc8rmxNaK5plr3Hk5IWdKFwWbWq9Hl0o2FRDwKCkKfqI5fbF8b1YghhQM+MQY46kFXH
nl3XEqPR5ZWX8En9w3EhyApOz3YXyyO6gNaYAQmWGNTeFDTx2hqBjqPONC904h8fbrnsY/pNfagl
IGgbTeMYlr7jsvvwqCpwf5iC6au1MbNMElw3VY3aZIp9f14aZ0SBcRvcoftpFqTfGz5U4Xjvtvyx
7Gc0lu43t5iycOoCGCFe0Mmien1OwlZQ50Op0EV6YPZIXH66RmVS4ikZfZP3L5QpI1EOPaFttk6l
3JKv6bMJ18tW33aeCfbRf3hBC97962G20bv6tbQd4ylhRoviqHM469FX7AcFXd0h4PGk+U+QzEF6
x7OHWEv1iZL6Jezl6y7ocThKTEsM0O5O+2K+A/fxHlDAopGHtdhfDbcNixD1edUFYZq328uu42QT
mjdTwCIlQapmtn4KrW6+LiMo5CoAtmTNZftq9Uget3EsI9kAjeMHjr00auLgEEd+03/65RX0l4qY
MWo3DlW7kUIKMpFOuBIrrI2ySPnn/8cdmszJ2xk4zISeamXck8LDYihJOcnjJnLwVRyNoKY7Nnm9
g4iqb4rFinDN6vOEzHXmlwfiuDpwSOhMckqycX3WsZKEjFLaNYkCOOoZ1aJWPuXQamwmZyNr6V/B
SfrHwqjqvNlLbFkjVb/+28Ib9MV7pxj31PaA/qvsJ2mscihwJCRWFsp2Dt9pcAIuoTKulBL+Q44S
Eg/51BaAP6bIdWl3ULN3lm8W1wroGNi3dmQDwrLsqeQjtB8lwHu7UpiVpQbKXRRyGNWEC0F9o4hv
Ox0kTtq6NHPezmJJMgLwN1s0OW3hMMkfL1NJKR+2F2ScxdtSRA8OCtU1cOXDJMZHj8aamK69aDVG
Vqj5909wD9mTvnzTpd4UHYqe3WqEPIQ93csgJj3LIADU2tHtiF0O6K9+T6wkjM2bZ+5sEjTqhQkU
AlKGqjXlihYkVtiV3R4z2W1aOeilIYTGa2EvJQCdVS095yH2fiZrEgER7BxyK8DiZvdUhEH5A/uQ
FzSdja8RvAqLJDmLtcIYz1hw6Yc3yVB0dvZaM1YxTjsYCBy9qscP4FZBcFMijogktsb4zwcOKck0
TONXn7L33Sgi1NIINkFqhwnE1XCV6aNhY3Gt75A0/auyXkrAKG/5VDS5WZRXyirDQNmfVzKcXQrO
F6rb0F4jLu+jOzj5S9FB4dKpGQbvAlrtTZGMsoWnwFFddkkx2tPF3EKD1/fTNNR3uFMVxDRhLNLs
vIOonpC3iKHr7yuEiIVORnYykhL/y6zREWPXEQ6J0IOCm8svWpXzaITMw3VylmSTQ/9atD2cP4vl
SWXoh0dMnNHkeMe+IQfiacU4k3J/SzirnhkIdcn6NE3rpwPlsb3uSipguqiqaBOcAgacYIosEFoi
bswaYyPO9Ngh+Z0fcUZwrwc+VlKaRQVR9AnPUn9m6z8CsIcFApks8YcqRYwscIwgsxigXCUK9vfq
xJhK60ulriRlN1oywvUNacmRMEybL0V+tEipc13VBMpD5B4rLagk1p850DikS0aQIlg6WCZvgadF
Dx6N8jv6VNgUaziTldoFIiVU54PxuuiOYeI+OZ4DhBgaxuLXpo4lGBlIzozXjMr9aHrlV8/6Hjuj
xiW49mTd6Gr3NTSZgFT4Hw+8vduZq0WOdEjxbrTADUSe8xjaFDvLKXZQSXgin6NksABD4q0xFOqw
gJ33NcthrC3uPchYnQOSRfi34Zz79zyksGAaqAG3wEeyalCZbRBqrVN/pPOmBM/qyC1ZaTN3d6ge
6W8m2d0PiSAAb2adewQsET7fLi9bRlTf/1QkZpZ6XRBlk/69Sulr56XICH8iHxM6QESKgEEoBT+G
09TqGROrSIwaxf8e/viKAmWWN5NDZJY+H1RprRwEVvGdNhYK8ZnHMN7rwcqXfcsu13gJlCbvuy0u
Li5GWlzu6DZAgClESwUoDrBlTORnAkWr9LwGb5TN7w/zzNMKxYewF8KdiFlDgA+BA7XDt99y6qMl
GS7+6frkGoPB+nOTk0hWYxAyAzaoV9/v0uq+NFLSng3CFWSTVwOujNwjx9KS77jZKmeiheeseBmQ
Jhfl8FPW+YJR4bCDsVz04aKWOOMEw3g98nOMDuflrBOZqhf7SB7HFRTIX2Fz7sWywXGxGhPtIJHF
Z9/A/TFJUlPd59KQfWG6EJkEWwk4uiJP+hhLhICF/ndJcpN3atRQqc9e3RubLqGZfqtuGECGwFMv
+CvpOtskBS6z621hngCVccnyFnW59DBhjROaNCpP04LyGzFLULMgjMEckh5SelMkQmZO4J9DkeHa
ufm+5J//igYF0zin3lMd5tXH74bwVQ8yttqXaA2d9t1C301gbNRjHbJtkgy76ttYGbTXlrgaoR/o
1/n6uvFtqWUB0Dickbjzvcn7pXOH37ObI6sXsbb+nGCIrAIJPTgo4bxpTB92x3w6IqnlHMtuUJEi
iOPJ8fjKKVl6XDiob2U49CDDbCvjW+Tpjl4lJX/c0r/scQsaGG5EnhcY92bvUTwDs8TybBzqRvvL
pbNLvdrY7S1NN/lAANDtXfZZEYYQ7R1aWlxTpkNGb1ybYn8h/3YAVHT58HqbjOfHfO1hLQe22zqX
ZnW9AD4MAJytC6+egb2ScuerSFH8n/ToQjT1pdRbakrQDOQF+D7GVJ1DTZhjIVIQXgnMZCu9KP5b
ONKmK+oBOrNiO/r2Q/7UslWv8DVo5VlusdtLURq/ym/OOg8OtkYTtxWp37VPjrZpR7rKYnug/30o
ALztcRNZSIuGyel5Ux0pmQV35snJAwjxRPflLtWBUdTUUf/AvpqpKy10uG6klcWZxV/6j5CQ5ZSg
o/qFAMpXoQt3+HvDpKV3sHXmTPRhHjE169Dh9Tq7Ns0L8TpOoJTTAaiG5/L7fmI2UfXLz2ZKmNzf
2p8PKtxiviLFle23kivbb50WvXtmEieHZm9T/MpmlJpBbiT1v4JV0jj0IIFlldodCKYZ429CCcOH
qqjsRg4XChRqudHwMK56hEPFB0ywO/p19cVSPbR45OtrU8+2PC5wnMS/UYq5ftLyeMJWHS+AVwpf
OkRzftLqqcUMNHENaZLSJ/3tUoAVBO31UllXvBhKfGBFBlWALf9e+F7FBI5fDs2ndCCN3qMilGbl
X+qRxG7+lgM8R0vJQv6aD3FkWrQOT43HH0kQEafJq3kjRjxzyWM/meWjQCox6RprJ2u0JL0b/oo4
GP1tTUSCyxvd7gMJyNlqdcAbTnjEMDLhFzcIVXPqab96P+LTCOKK9EU+D/B5OGbV7GwlxItv08lS
+DWEltI1JnsJ+Z6v2e6QkX8lXvUjSNjdnyUc5BiXdLJ067+pecw9XdChzp2NVXs4ZB/V1wqJh7/N
ZEe2qe31+H1RDtQFWeAr7fH6/WDZRw57yKa0SnvjC0nrfsBKw1i4asrDLWy53Wi/iv3Z4W5dStlR
kRzHEru0GADHcrgzw2TAcbXMg/tkDNJ38e9JUznE+qUgls9kNIpkLdzXRNFctqMGQTKaQJdUvzB7
W7aUUGRbGXuvJ1N3QdZzk5rFXERJrnAq/ffVRjwSlDmVoGwI0C7JS7pKMgsQuejMm+47u5BEx3Yd
8p+bW7Qh/sJ3pxqTSdjPgNTOBKoqirC08rGUJ0FFI2mgvlWlgkHYSeUTRzbGM2hAcOTzx5Fe5a/e
yUI0sQ0WpX3m88CpOQaNovSYx27H310tH6bdR1RYPF6qRnA0VBUe+uyslW4nHtP0ggeAOGJlul08
CkoOd0QyC5uIZo7p60sDTXSXVcnRvDXrqTeSQiir037U7VsImWKvJWQ1ZT7gwds56YStPJuiBCfo
5altgXeadLdtelYuJVLnhxOpS3ZFICFwe6rOtIZqnyKl5fncce4RmbTul7vCiTstDmjmHr7AQb7/
73/m3Sbi24pM+vSxioCHWv40cp6VLnG0LZrQyj46Vum3l4v/NBEo2fVintNaA3BFEJvtssOSdPW7
GmZo9qZuXdhmqPpW/51cf6llUEt3n6YwTFb+GCe7ZjRadXhFj6qYdDxXRqqviTYVIuUwUX5Q4ifv
IlL5BiFow1PbKhWGPFnd/+nVpZM0LTKTgZvUP40vopw99cwqPhXgmlhbD2eGq+cn5Q5KDfxDOMxH
Au8MajXJmt2JUPA/mtIvkc9Ybj9M0GihOsOPxrc74vMYsWdOZlxKQsGRXlWA5CeiHbISfMdDsVAV
wb6+XeCH+09DSjZ+EG7ZvlngYVtJhjinj4UI2jg8x554qzO5ThugW0UNx7PYMst3SNCihaNjs/8Q
vrkceahRCKS6hilRYjJu5HWJ9tBvNo9UDdsXz/wEkpt/DxRCFANFsRjk+OamJMqMN9IUU4F+KaV1
2Glg+qD8VE75jenMSpTUIVFanaIS7dRK/3sZ6/FV1S9rOS80/7CBkScF3MtbCaMOnXNJEjwLi0iB
Z53PHztoFJYFdK6RXBXHeytJwcTvaTQnu0Jyd6wLWubDWZ+U4ONI/T4m9PHZ3JLBNc5Ou1Vcr10i
4C2ys1CHJSGAReU+coxYHzwfMOge6TsCU5WTc8OH4yzhdywRC/cciHP6jCwjvco3MNsgRttJZRvd
nZ6S4zKbbfsb5IUbklwhAlz3kEUBjI3B0hAkSq/4fAgJ1eBrwT1zTHCLJ2mwxV5MXElNVTPOyS13
6i9JI4BJzqHGWTi011t6ApGwStVofhdFVpKpx/L3QP7qe6IBZhGiH9j77m8Y014TTVXUA8cakR26
I8/+FkUh2kVEJZei2l4qLEoPpsAWa3DK/R2d6peMqPNON6PKTMo23sGHdVKXmKha7PMqJnRb93To
HCYzWhHJxrKywalySsFjGNBxOfeSAxztyOu8D7l8lKPz8FPimcMerY1xFvwY3eyBJeeBnrarq9R5
2llfWP7ohn18GfYkkSTdXhoMNzkM3Mu1ZsKSz9uHF5IXce0s+IGhiAfTTyRIYGQmTPZ3zf92Y/Tc
4eeUxfVEZMUtxjlrHToaSENsxBNWLYG1153Qf37ftAa35u3cLy11jeAYG2t0RDwqtUTg5qlakCMf
I+SFRgDbOpn1vLeMP2OCJCcBafAqVvfjzsle+jDvnBoThUo697/wAjJ2y0DeCKzrC1K0VqAf3cCv
x2dkacAzBzimHNZxAoKvmteldXxF0hIqiK9FZ4n+s5Bmx5QohwOYGlaB3BT9SEFKMU+8nAyHx8XM
A1qjjoobnSdCcWZnbvRxfqGDfGZT4ea3Xe/tdOdIEjtc3XbRJQKs5DoRofnePnWvHIZTb+75fRkn
i5C0Iso2ED0I67ONl38OIa+F6bOvICvL0SzPFNJa6MoR+qC5mbMvPYoOU1WkKRwmq54iiDymBa2L
MtXqb2IEReNCeEX6ckEv56CrgQvH1/EBCD9pbEURo/gqXRHQVNcoW6H/dPHsFR+fePwZOhn7RvuT
4e188bMrXiBFP50Hq7tFWTJ42FHR0QKrou95ESGw9mcGoZDNblnJOFguwDkvFCuNoAmYJs/r20ZF
CyY0/JLjq4K7Fjd4ceZEglrfqxQzEBD6ZBHjWJP+E56GcruB9JU9GBO6yArkDaeAv7i+2+GADGg4
q68GxtQ/T9DM2D2am6GB6SAFFoXqhuq5+K+7WEN/i6iXlZh18WdszQ31AGfhS3zO3uK07eZ75zs7
bKsSQ9UpdqzgjolsgCnREhWWfwaxTmAMngt5kpJDh7RNtBLr0oxJ0DhonxOH9mU8d2iTG0gmzqE6
zG5fYCS6wQ7Itt27kVmuUHdA6o+YL+hKyeQFjAAWkrkxnAwQhONU9nS2yz3BDPyvIwVS0/t8sB1X
OZTepeAfPscPt8UZxN3/rvefAs+ZqxmAukGpqFJ0jXnpzezyXFl1z55gmZyLFExYkj1NHY6kcfeX
PD+76aoOzuB4G0o7OHxpSeXHuLNZH3ovqPDbywxCOfO9FmUgkSQShM4sAwTe12E57L9Phx1ORLgT
CQbXig7NrWf9K54VXMfI03jfmrT3vYd+TTI7MYOy4T8psUkqQ3IR1ZMpXHTqcxmwNyGe2ig858L/
wwHi7zyHnCiKBHj/jDnvktTuZpciAhQjIBmmCCa/DM0U7Cf/S9z2kmcIw8xd+7fllo0aTtX3IcCa
zX4OqL21cSFhGb4IBWEx0gXGU5mERQXEQt425R/3Mr3GpnK9KsrvnsTuaq89x/F/1GuGPPB7QBFW
qFWtrCn93KrGgbDnJLvw35+rPEjwZfB3EwKKxnTK5558iP2km6cjIu2HwyY4k8c4trGPMNjCoVcP
lcYyjXWHdhgc3uvdnyvUl2vAGBjg3j4JQKBT6IaWwJqgbSsIaJ91v/PubBdzgf/Ym2Md+UQPyCrY
6JAu1cetfgPau/1d8mcAWIgvK78UZs3oOZflpiuQNwxNZ3rhcdoK0eIOr3uh7kaeSaW3oc5xz6DR
9H+9lzFgLe8uFibnD8N/foKcTp5G/48IuQwFH6V5OU6KSb9xNNh1uOAnlIU37nPlWuURu0UXCNn9
kpBqCc/A67eIQckujq0nG47jV1DCmTXJSbTvKQc/dJCVXpwxtlFiCW/TXaT/YXl39xsRCT1Q1/HN
hUkWq+4jk4He+gkl6T/c8eaetjU5Nvm+fqdB9IqDh7aJJFOCRxROCRpIPHldYpNAnXWtrx6D8NE4
vmzmpMviFS/9NwlYEsgO6ta4tYm1QQJpimgiDvD5QFQstgAbJq4PnycJvy9gXPW6gdDRfIoVdtuM
TGTIBenn6ZEUrrveFQIVZDx60ZHASjE/PVgQe+lANe6dIQMC7UWvR/sVWAxMFuIuMcXWqrvfpb9g
67BZDiyyiL/bk0QFS1jHX2BPHoGxGPrEQBx8u237RUhYTGDWwYsyQs5hJVVq7KJJ/bLU3gPNakWi
uDIkPyab6WVQSylI6lisF3Olnc7BTmTGtzM4f7B7KU+j7sOIp5zHGQh36K5JRZVJrYCm6nuSR2kO
pFX7JSs659yD2zxJcyeEYhxdTixgsp3uFAZR1rRAEzbj4vQpzen8NTFngWVujDXVIMp+CnybS1Ot
8ar6Owip6T9ivRALiZyvAHw+E1klBqRpA+As3l/IFcyfIUi3xiilw9R88gYkONxJayU5xUPg4oiY
v7og7dogdDSCmTaQYDcKmG47r119Nzc1XmtVo9YAULW8pxJL8xkP6fCBBZ95wE1WoGuhicnQU7Z1
p6q4wijAnSaUv71GHT7o5N9TjRWQohLGu2/vI1AiGyuMNVeafpUpoP2aLS0Qi6inX33gbBiT3XOY
VbTRbxhNeAoJhZC0qUNvI2tDot/ZQIyrnsSvBPiJG4HSBWm8TXF8J9ty8/iK1jeu27WuuzWXsVLD
fhuDA3OFA/UwMPTMKlPeyamsPqjVQQGpd4NolWjQ00SXUNLe5Q/GzQkc2fNBVKjguQSH8WDTFnoj
9ASbERRk7SBQuZ1fqHo8aveT6zbCn+h7TcXJW0wq8ng1/kmgZbSufvfTgTdOTDHQL0m6KluolkNA
0bjG8EAj03aBAoh7Dwm8jKWpgLXr3yWmNLgdbgy/gfKpQ6Ku1dcChxm41c2K386VkYR5IDaac+ps
qOOBAb2sNHSPOUn/ZfeTUeLIM/grK+V2s+3zrhOTGpTmH58agPDKekoEHItIj647TEdN9DGCymqq
10CWVLrzQ5GqXsr38kBLhtlm8V/C6uk44lyTjwP/vJX90LsmGYoAaBM1jbYBEHyLsq2nh6aHSd1W
fVkCh1nYDPykNZfruktPfaQtrCxR52vp2S+fkITUlfcHsGXuHfcJlVYrgxsEGhttGCNpQqZpwdVo
SA65NNVdTuUue5bev85cgaBK8l33D09bt6KYHLx52VNMOCIcgIjefoAvWhCdUnWMKht8Nn30u3ee
/2tvxMwwPw57kv0BND2SLsPgv6oqnwmkiKgMhb/pYIlU7jdr51RYs00T7DDmKyItTh+SqxAKgEa7
geRK8ERTwbJmPwsmCs4EWaMzp3GdXbKZ4bGZRiPhR7O/fkynAW6c2tw3ZcarBGG22ONKfctKYfna
3iNuJfMhs/yYaxMzXgnt2yM+WaK14RBEYtFZantY+oVqyfvAwVIct7oO8zsH+5XZnCYmYJO1WoPy
fM8liOinIgs95BGkxVA59gFqT3ps6cRcIti3i7/AfMwHtRppVVwTtFe4CaqlKgstkgI01TOK6UQV
1J3dwf+Xw/jRqgww/urUGvUmAWNBfpIFDTBlpJHKHZY0UI6+uFZA8QgjJ2LDj7cZt3JpcY5i/WiX
dUd90m0blaIpB3cAu5Cy8f4C0SIoyYrmfcAwVYOcIK1A0xs8rnGlfvG2PSPJgi4Qz0D1UOj4UkXw
kQNW1S8hbRZ46RwXUceXvx9PMOHPaR5C7WHdj+55XlBVCjuh6k6zGyHVl+Lsdc62VVYz/sP2oBIU
nnNCnrvEsDxSzMFDFqAdt1rWTVLLhRBBiim0NvnXgIT2xu/Ej0dT8qL1UPGdaP8q1aPh6XP2a8F8
RBNDGcnCTdRgM75baWP2ObO4T1VN4JFR55aVTuiPYi+zpf6KfHgaTDPegRsr/YTTj8G3NscaPYNY
s5BjGjdAji6MOEisNjrceYzyKu0WliH0idihEZLv+Ehs+JDqfoXkE1PukfuJGB2n3q0Xo8af//bB
M+LhlTYyz4euDGQQAJ/HrI70wUf4mi9zuMk7Z2c12xWKRzkQSiB7901s9iy/pcW/qo+bC1HnYEV8
pOcYySORuZZ4ERveougWTBUKQOtx2eXG9NXtDh+sAjBm1Oxgh0/6wSKrdQNN39+CO+MUOtdd3AzJ
Ej0E7BtxEaabkTjMkWZrgwYw/oaZMgUD6g2yweFiRDhOq6WAhBvMfB+AIdgudx640V2QcTInZ5Vf
BfPOgu8/g4DA9+trP39d5cyp1Podj+87stFXJTx6mbm0uxoHgcLf6DLheLslvR6zS5vQoOwgf5BF
FaNElGgRfkrJv67M8roABu+DPRs/xmWQblZFrb459MupeYkqG3w7UZhccD6sMwfFaRVW30MWflyy
nXG2wc+zZvvQ5iU22WllGB29QAcO7FKQjt2ICQX62UCbFOWf3RYlEXIJiD4DjfW80HhUwDsJCLgj
jTEQDalin73Kd6CUSai1vT92t/yfXHT7g4j1GHFuYc3doo7uwiMfWLIOx0LFcvqSvE8VJfaVrR5P
JWS9dwHqR5r08a03nfDCFlfM5Q0KPQrDbMFPRl2esJQCr5Bue5bNz/dyv/J/zDmLyqlzaQMlZ2fx
nsS0qEhBUlk/IuaHZZaIVsbbnae8wFBenBr3qyVP9+okecZIMdc6O4TsDBUFeZirXNrhLNF1Tqvz
e4Yz0f+wY0YfHRlrHas2ESBOwk+BVQnR+LPZ4PnLApiVg1snGjsL2zouUxJDrCE940RqB4EVPDT+
LC0hrhZ+2uGd4r8z3DDgGFvsJCrblSyGX10xL8J5t1bTrKSf3qryrRiPSBukObOECHhmdo259agP
ZAyh5OeZrnOSqEqGOVHHvhWQPo2MMT4HMXt5bJ2FZ4bkEwPBnpTobVo2Xj3As1RfQuzmhPdfMxBT
zhdG2BOCIGhFUEKA4wTSaKPPzDco4cfPyLdUGmkHVj8ztcGyje2P/1YgraGbZJCEaG4lZ1lpXszg
vV/CuzeDOqm8oSH2RFz+NvCWx4qJ69rgufh0E2E1P9Fqz0Ht3caK8H0HM2JEFh7ysi8BWuVMGc6O
kDUdKM1fY5p9wO7X8TiZX35LXXtTlppchjJNp+5iwSWdhevsIFD1ZMiN3h0ABCRjVDBDnSljaH0j
481/xWfCJae35WvBK7cpsL4BD3fATsiY7rqYZzf6C57FP5X5Lf34EMrBOSAScMK5+KLT5RouaIC2
MjTCkDJmlNmqk2T+Vq9W7AsbNGpXQ8lVGWKFeBqLXblTQfT3YfV0vyul1roN5V8UKDm8gNBhprUJ
J9B3GezMgyHlNEX/m00r6l1xlpNt1pEj4aY2Nb6T7IxrtG/9fX6BxLlDuqTEbDx9WbLG/DSH1e3M
EXP67lCvv9kUPGVF5Zub5lfCeKmXm+yEZ42ueYX9FUaPjXEwwj36XaPeFpXo03STSKdEWGg1SPmy
Pf7LkBixxvvBCdorw4ILkgDsWuPppOtmW6OpeTItu8rVPK8pJuJ4fplygMPo94u2hiJ3G703EAyk
22LVGEDNhrPwdW5Rb5GgK1bR6TYIIWkSvmNEQPd9mKS7AVflPrue8q0MUTOrjNjUTGHQUk/a7Iws
SFowb9gln2SCbakgd5R1QGL7+gCligbvZlfyzOkeVS+Km4VW9bH0ZL/hKJ5WzsSOzsME4kS2GY4d
miXvcub1V5fuMi019deOL+/s7c4RXEH5aCoyl0YtZhEHH609/XcqaHTghGXxVGtVpmu6eNKjbfmW
QgUDUVytc9OWU4JKD+nCUsLxCitpk8cNe9S+BOI5LozyjgG1tMO6AO17O4qUyXHzRpkyn6WuGbGy
u+d/m4JM1ovMTuu2bB696hw50GoFnWl6oapKE1n7yYxULQJ1EfrPlTY2JNQQitDf8CtdlCI5BeE6
wRuhWlZcuwptMIy3/qk+yLaoWDuzR4PbvTgJuQ9fjifs9/VOL32gxAOE7gbSjEl3end3Y9cDK12S
L1exAFfha9Go0c5wJy9fByj8t1nS94f3Jjm1IpitgHxOgR32+nTJZW7xCbe+XTMxBrfk1D53Qusc
hE02Wc1He4Z8F7ldszg/DT1BB+xMPj6ieeAZtXsvjMyk/BYJpmIdh1ggEAVnhqDQICXxCEBeNhlX
86k20lJtx7Kyav1ri1XgxUWK8zuwU/UJxMcDA226WAkJ+p2s4E+Kzwms7x2M85eUJWzwY/Ph1jXT
6gfD86R+/2aMqC7sHm9y1oGVwf2M4diSetNoy4DR1MD8TmwqflsnfbZSMD1ianUpmz2cRSswuBd9
vP966kb8Cd6F/KC8z7uud24rLWlwnSdFJZByaIxfN12jJ8YZ3XstxDO7jucCufOPWBEnf+sr1Rpd
E/NTSwSTEhqwX6Ds3KITn2oTk8IT1lq3oQ/MmFWH9jvO4SSJAvi8LWluuvEnPxyG83gublrF1nCH
D38BSHDsoaRmApMYeYbi9GbFz+UhWSZNZFuIPd1iMVXcCYOkiIqdUtRzV+X0exhWdMhyKY+l7OAt
mSyjTZM3hddFHcC0VmvnWtfHi8OT+/QPdc5I/lQcb9iGIVx7gXnTRd2gDJ6Po5+TzKXCfJ7GO7g2
Tkz968vgMODOXjy340wk6OkMFM0paG9LpWsHrjrDu4eGdwu3uwMDIQG9mkBBNOtkT8EjfrE/hsRS
DJPwvxrDWuRyNLJplBwNpsfj+vF/Qu19k+avRkNCa5qLNM96K+VcrXDS7Qt0Q8cyQsuf6vH06B8g
B4vbmPZI8KOL56RKSyJ0BRxIeH+Px0iodMvFMatg90CsK/oBrdApX5/h7kmYORrLhTqGg6H37skp
vIa/qtJs2gLbJgMlV4v7hrbrcUHGhPUr8TzTJR8LTUKSy+KEPHU/HBOvcvV6n6geBvkzE4d0kQK5
UzvuoIOCxZfyrbsxiLISx9rUXeo/f+o+iseaJsGkKvQm0D0Fb7KlzHODVYBODww0amv3nJ5dDY+t
5f5amBj+u2EvVd+m4HQ/D6TgUxjZ08Uv4THF2uob/CzdI+OwkS3i95scfchVjDjk/r/J0wKBj2O+
zH+k7eKHtMXIf0JUFSTqj1mthFuzDHTV5CY6/rFRDkS3Xa2aDWL6HfE8lphD+Cj/r0XRN8JO+ySF
/2b0JmcWNXLrmRN1D5PcG1jZhqWjaWYX/2MpAsI78q83OAUSlzpZsIVag/bVRBEKFQpRY/rqoF7L
w9pRjc1hoHKtEZdoF4Vr72MaVpDx4yrV98U5uYMo6qN+YcQmFwbOYLxbfRo4unuKijKD1f8HkqJi
colRnTfGBYNV5HdRpyuznXA0zlYYq+IjtUQoBtN3eTr/WzDwsNHerfZDZfeFwb6KT19fzwDdBquH
Gc7SFd89i34CgfDv5Qe2UriUDUR5ckh8XaqMJJQfRIZtyfFLDFcSmo3W1Ilo4nliqPHZHrWGSx4d
HQ4A1URPuTxhdEWsjTuV1Cxx5Ylgegg0QX06SySZqbhPQ2sBdcFVXouQIbN/lcia3fiTcNpxcHUJ
2Px62DVpoXajFRlEDZmr1T3axhhGohkJrFpHFvMIHHGkTvTEEZ6u2Xu+UV5fTAFVKcamkihxgsPM
hYU2LMDVuP/gjZjXhbpa9yjhvYtcfhq8WQZCyLEb1a0GrzDWeMG+SMukty+z9cobUqP+tn/7h/am
pi5kM1spQer4lgtzvB5eS7msczRnKJH1otT9SJrei5foI5rLfWeOgzcV3DFSNysILn36iSWwWJig
e+ZqDKtsnnKDjpEmVeMu+uToTkeRukkOR+Sa52BU2Gw5ENWGqtxM3/DIfPM8uMpVLxwp766hAnhc
GkIn7xouOxsZ1ce7GN7ViymBL5IQESZwP+hQ+RZp+3W5M/tsbUfroFvNMAqyNbphYlIgiCfeZRaD
h7n3y784/4cTlhNReoMnTTsu9BeSEnR5QK9sJ/J3cIStuaABQ+y3Qt/Nt2IfDY1ZL8MuASECqHnd
680MltSAwJEn2OYHsH6wvzMijrs6Mv630jqu17XPlsn+5Jp1OnUPna37/wm3TUPtX2zBUZ39Fo7z
aRPKPrUB7WEQpbBs3VCSQjzc0SENJRGPryvkVkrZx8KHvCsWup8kL4lgotSmgVTO03eU3qedVdmB
yDhZJY7bkziw1mZXJv+1oCEeLot5VkLWNkOGvKpEFRzxVskUJnz/+92PqONbsIW5bPeW5DoqbyMO
bAuZZSp3q6o3IzZFLRDHgwd27CUNNsyaReRu9SMGDGc3iYDeYIc2LaGevvLpuYpfvLD3v25WnSSF
62YHgnNzNjIGPg3xSoQrOvO5iC9AfoLaU9qDdL1M9z6qmN3y6hZhVHS8b2t5L+YtUlKezKDZl8YU
JcDkbKvNLULIzqVdsBRVA5C1ioLBwt2XWghVkzjXBal7KwNmaVOfrjUG/Z9wWHlXQXg100Vuj4BG
aXKy4IDpsVB3R3BOvyZjH15tH90sQRQ7DV3v1p8kKe2aNDPPl9LiACVe8UVMKq2hKfBnDdQMIRwV
br2cVM8oOX2gag8vcMBx5p7EPLR+rc8/pRQPmvqMe02dvXbxtE5s0wjWYEg492MYAlYqHXp1ZeUC
hdC47qHV5vLRO11S5b2BZGiFtLbpb880dqEIy5XMsuAZXX31LhJno77BwwrC15E4iDWaxg8Z5OR0
24RBV6AI1XYLcm0I6HmOdu4l2V9HBY2dy5U9/nkfUYYr7J09YKWct1A4juV9f1Jsm6vTpVZEZDo9
7fG6+HqBCy6+YjVU/bHIhnozKnCTLmpjQEoHp6GbjGs+VekDj2keP9cfhVSsuDkc9TuczirIl9mn
rj25gmwR46uJ4cE+t5/4rVknCoCgT8w+vBTQlHCCCqT+t9KUhq5bIYTM3OiLICduAPvD+iZY6x7F
iOc3UkiyBePGk7cFKoVdgMnNEo3aFErVW50NOlBzBHTRAiO304oAGBtcFcm01ThP0td/7nFBVkNA
eRoHdHZfjgSBfd7YkddX3ORLC8LXjJvkeb/IPNrveHC+LM0dPO9T6GOn4wgZkQ0en+gsJgSkjBJ3
ruAcsoX6Syn6xUMKdoknUKoN/88kWEQbL+73tqQsRuPS3w/jswF0ruNymtdSbxSjs44ldMA5DjML
S82f3msAIIhdarov56lOTJWubU7lKI1x7fT7ArGXVdvRv/kZPL3nabfRoAaHSP/lI9GHERhlmOHY
dQ7oWVjwl5fp79WxDLKTcd118FEAi//c+v/kSURoxaWuiaMBPjJF8akqKZo+QEraSVvG0aKwRGbO
rDQLuJlOou+A6sCuhmpvAUnBI4aiW+KQM2xBeffVHCU9S9lZa+2DhTxevZ6FtmM0otGxIZ0c2ogJ
49wpDKQlEzGplPwWiNa+pOHIWyHQ2apgA0PyfBGIDzzKpK1XYjf4sFnxjTYP5O/noqhCwfgHoFmu
8lKrHtKZGviRYYSUKxb30lSeqABcswfYAGw2U2naOwIzgwD4h8pbLuH4Wt3BOvDKB1WDMD+eECJD
GCVnV3NwVK4iS33u5QCZg1p/UfWb/OE5xmOyglqSLhYXmowcJoGobVM3f8fC6IWhxAHYIwfTDDYu
FuI5RA5o5sWcHSOz0Ks31k9YIdDUtK390u13Tp45xeOk0VP25e/OvQ16Sbnr22YkBSry8fxeYjoc
ioTw8FeLiuzqDITAtEhYbZvKB26lTHYgW/0ii6j/AIH/+Qc6g2a5z986Uf5YeuQRLoFeT8WJsIQ8
cBAnPConPFI+voA4y8j3krwu+r8pITqdPLmIkhWGkR/+BD4zUKl72MyTL+dyhGMNH2dRogZsLY+U
T0JZt0xXEcfrXoPu+Y8HP/uQD5dGfOPrDjdW5BVew5CzetUWU+aG4Pd0wPDqUJUvvLH8RKI3UePE
bCBSt7fcy1FOYla66gi3ylFrehZjU8EJSDejEMsdLvsyeQ7QY0eJiorAeRK7KyoCktC8ZDgMkn9j
ARdIqYEZ3ICne9mIQuV579zflP0+sqAN25nuGSpOEPzL3KvWc+mOMacl9eLbqF88sBgCglShxCFg
ZZNw3fB4hiExLQozqFeUWXZhMm3DIfoPQyMITynEhD8ombAtK4z7rgVfvvKlM0a2AOv0mtPHY6Ik
Ex7dmUKpWWYeCDaF8mrpmKK0EMmau/QNqX9+az8BKmQsRE/B8/VwI5+pvZIV2YwJdMrkGRLAgZc6
iqtihuD6evEvC+mLteazeXXKjGagEM2UV9W5RXmVMiypEIiVbQQxGLaYIGr8j7lYAG/yb7X5abgb
VCiFRVt+19hFIwLZDbCwsQV7B9lL/zqX9aXlzFk6Xv9Ui9XXjfN8I97ooSDN+McMFRtMSkCmOT66
mE6dvrvjpqDbbAbQK6JweMZx18jQIgBBeuMIIGypJLDbTGSWiiYfBdjSLmeF/N3MeFAfzYJYXiJB
nR9jRb2i0umb+yp05b4K5+LXAtfb9S9tW9U23jdZN0qGRBBE6GXzraocCWqkDcnNfh0jQ813S/fA
0mWcQ1k1khh2mnQp6k6Zn9MRWiw5u6XLET+4BZ+1yoPind/knePeh8k1ZmtuaGRANLvlpb3JqO1X
tU01nHuE2WcOf8PbGJN2NuTB8MeCmNspu1zMbkBJTC+6b+SUUZuH8lEf+DQ5Mwz2k6+MUSFAGs+V
k1tFUddoUfwDXVKKarcj+rOourHvWZwN3fqLNjjKbgpSf7J3Y9K7WLE7ReB66CAofqRtxbgMlvSR
0tTR2v1r2xlxbECdgL51zbAkD1B6zcDjfb7r8HmUz2fCBA1cPCqJwp9+OvXHk32MevRPUHmd7Czf
5XNDS5n8jkukQvJTaesD6xx+MruAXesbxfeBckXHrlkmwIsDiL38KOn27zRAqbEyeIxOlpvRwdL6
72wZPEh3b0I2/GJTaLBvK9H125OVEmRNXSIwNlKvKXE3pJPGbJ1Yp530OCoDEwa7b7wtvtkjHpIh
3Um8ecPny0kf5Bho5amStyok42cihbjZELnCn9lq2XVbm5Sx+IA7R8XWxRaG1diIOj3L4xwjNvF/
AzYT6dYUi29m4MM0JsXt5H0RC8g6lPaJUTJPf/r4Pab8/df210GdWcHqdcY41CmQpqvTCXWESWKo
vBQ5hXkABCX3DMITJfAy51Agxz8c+iN3oineRxwCXEfcjgz8OUYa75CT+oskJAGTQyeSgIubVr9G
096lTt/4iVTfyyZHLeUM5BqI+YyiX+iUk4ft6y1d54W54zH4D5lqHbl5bOpl//haUTa+anGc3Vm9
qgFpuiP3KSdiXsBX+TAIxa5rEC+70wqPaZvlsYTDG/vTHMVABlp0o1oo+Ird4GIT7deQ5AcTQL7g
tqUC9LNT3L3AxgymvydIaZorvX8UDNcZLeUKyiqpTA3EfcKJkvxJCWFlNge6S8PB/RS3kBXJvPjF
qi/GEDe0q1Kwn/wr3bmgpfgKvFldqhoDULTSn1sSx1tP7mu2i0Fg6G1NhQeRsJVXeyix/7TVcE3W
nwz1DOCjrFr80kBBNVNnMIqFHnVviKxNdab+HtZBrLSAohqjelC/P4ZSZ8qEsG3xSDeODUPYl+Nz
Hn2u2cpzfJ2n3wQ3ZWNX0nHRYY4K5nJFHe/s0i+HoSQ/xBEV0WyyhNPB8VkfWo+TxSjJA9PZKkE3
Xty9RpEyiBncihWmUrUHnjd0PfYcasfHmy+KfwJRUXH8TMV4UpRFpuUvU3CCMugBCGE+1PYVuXNy
pmQOJGhgHd9/Ta7DI69CtEtZhY7f4faBsy2wUXZesgy70PHXTfgRCmWLmcTYKQhMkGMDN2DFBLQx
qtftbw1qol4dLrX6WaHGlzUMfG998ppNCfqv+kzKfbQAHxss4cd8dza8wkKSwNOw9PdeBQrECsll
X9hhkA7DtZD6kvQWD6FYinXAepsX9QvR0Y5uHRKGlzHUTO4cxoAZueMWDWBIMvBrB12Cwq4xusY3
tU3MkXH9K4BJa7N2MhIy23NgZGjYVifWaEm8hW0wlwkEq6WEj+OkfNzT2v5eXBpXZEIGAkTQR8bR
9xZ4IemHIs9oN9liByIQTwJI0YZoeXMVYuujJJGNrS8X32oN+d4+CuCc0SwoTWDQiQdCd4BMgbkD
VIiihfckpCmn9Z5+ZxvdiLys5z8LcBXuTkYMi+ix1+f3lMLGOKVwjAvmDwOKkpz7pVIIhwGa+OxV
9wz1EzqbaZWuX9UXGP6L+v7/cscrjxVzJpY7w2bC0NUBgHonWdj4hi/CktTG/BZn8sf7azEP/pTO
D/CPmYDg5EVvHP/9kxFW4/jyVygivQ+NrVYwCjhkA3pJ755d75Lx693HbUYHUJXval2Y1HToFQ2P
MuDykHf/8vlV6JQS3EZs3Cs53SxsD7LIx7cb5uBRL49FjInC8VFyJt4ffarsQJc/7Crr/tKUwLzb
LeNLIpjsArQB+8SpOJalDZhLADFAqHpwAayG09FRVI0VJi4loPKZddvThk0wQid5w3rnnf2DpHQs
hDCL2fWJNZb7yKlh/92HbpuSAq2aH8a4mhUAGKDe9zz+iRVlZiszRcoYsB9tQp0xESNu4q42NSbp
0BBhVJg9TRc3ffPprBEG1V84lpUq3G0id7k4BnIJW7n/jTwYD+p2Evw1yaLpm58H05xMnZ/qYHGW
Y69swI8GgbVPdP5LOVFH6DoY5Mv/XLcGUwI0rEk+QXuV60xLDeSEQIPWtDhpJngrSX/ztvRa7O9N
zXj2GD/nDu4vV6iqbEkWRN1WJ3lxjlrw3xu9Av868uFP1a9Xum+DvXegx9mcywYdBxbsrPT8S3OK
G4Q/btf70WrUp1wNu/hwwfINSM06a1JNW7mzqTgPGYk2fF07zZ1hZP0la34pjr2OjTXLxrUSXvWs
Lzb7XKH+np9bWU52T7cxyz8Ftri11/mIVlQBKjebIU0q3ltPGsy4Ty66WDwcOCEmebTC8saOFQQR
Ny6LeU+MkwSmMObdoWB02telL2YbFshlol9/kZYYT2+iXH7h0kU/WuPJ7zycw7GecdIJG+MGSKbS
2Y7UjmwzZ7nGoMiEPPTnB50GBBfuMKdXGGPYAE5IIeD0XhZ9J/WBsC5Yy7OOLu3Wuqkrqar8EF1N
9uOVb6XFa7AwIhAIuWN03h66BAmIE/ksz7R3qdJb8fCqJRBf6xQMhp75eUgBeeUca1BuO9pOWZMm
XX80dpS+x+uCB2PKNpEwQ3FYGHVcSIN9lP8qJ1MJYN2KDh1gzGQqUCSL8H83IzBAX5L9x8gur3Uz
4IdSNJnneMBDwhVlUEIZHlfvX4pcBbShj1qRDAM1lmWZYJdySh2GH/Vdadlhx3gSzn2VCRNLrF/0
akI4sgTIZYrNp/BCgNVi9RWzuOSngNFuFj7edXpGEg/75GRjt0ZxZf3/qUD05oq7QangLq/Pv5dF
su5AT54GntIGo5QAVZRq5jauKjDu4aqK7DBQ/xfzc8ZRARXOw0apc796ABGlVP5jpYUJvvHsCJRj
WyQ4PVAWPigYFauCr+O25shXw2raOGm1hvSggUeH4qGxADZz0Y+DxObh/4SZB8V2qXYsoGEUaRG5
f8SR1j9Ep6iRdfBTEzW1RDfhMBqi5hQduncoXiMe+uLKkvPOf2WRSNoOBWQsW1xmwQ4ZHlKxYAOn
C+uvEfO74mqYhIv+6sq6BMGaG9ljUDrBW3avZRoW0eFN7b4c597hj/ngWUKLVjiRukj2rOgblAux
JTc+51K43rELcfbZu7oRwL/KZwYewQBNpj2XbnRJfYRht6KqYL9qTQf/dyCNnlAk9z+AKe8HDGpe
d7u92FktQ/113baNhZVHbUQKtnlbt2JA8YM6NyBsVvT/tJnWocuhuGEcoVGXfEJtVhDNza+/+IH4
8wRpSu9/G2PGFnBcuLv9sBiiQlQsNGP6XYBB+yCdKGwhr7dN86kpyM/y6PJ7mxryvbZaES4/j+K/
dp2+GM9m6vOQIz1AEfti+ugOWfsBrpvrDKWkxXi1h4kjAZGyuNRbjbuYKxqb+JKWGUNH/pWIaYFA
6JQeCvLs7ggTdHTyL/tjgRy2daj24AJAvNyBCporyXlGd5fcEPKsAIyYENJyUjyHDT5cMnmGZan8
dz/wYNvKYwi/Q5q+7GbHAF5tQ4pD0OorJJV7sQEbnkbUFaPBctAjQP5ak3Tzv8GlQa4yZ0iYEFjI
dfnJBHoS4RWH0Qh4aVceM+9/PYbZoEZZHpCotk7KExOpKSr20T8nFDfSqbHXYlR3SNTKetXxkJp6
XGnDCUDTVDAizdc4BGYQlL2Cnz/QnR1wURdv6Jz8yt1WtMFkQu+a+/pDbFthlnvFEtcY7yKxt2/1
EAPq2QEIepe8KWeuaem2LHPhWuDFWka4LGCz/l9dVC6E7DuWa3tCGT0edw/dDaXKauVPy+XVS7m5
iC3H8d3uSLG1EXvXxvhT1/RDMyJbSjdcyRfTEc4T9AuAuHu24oP/XKcjmTtkDH5+2+YAss75x5UV
r3LG/RTSwMO8uNGZvwVfhvu+In30OdD52RiYGogMI82MxirvwBiOtCEL0FFZO7EIVbBRnIe3S6mG
FDIE83J1XrO6t4k6paKqEMPLl8LguEcCOiK04F6eb0wvFIeWUH3R8ZzU84DMYYwjKhl79JyLV12S
uXCdz0RBuU9HqYcc3tO/3yVkcdVmV1ZwUobr4gC5hnmwQd5MCBbhZv6JrhuFk4/7NzGcWR+l9CcY
PbtcoRFv7780YQ308EYsIsioPx+hDLZjQ0grYKlwqyoJhJDwNziT45J0Y+BxurZJ8gLdMba40AqT
vygtCFbShIYkT975VFC6xPkOlXo3hh8HFFFG/IXebAkVsjXNS03pQO2G70yAK4zZGEjq8HHHQV7w
Lgmh+TZzHfbAc/tvlBJoMTDWE2q1NCwnhda/MqZKncaXuL8XxFweUCcJJwci36CSkXwPqAkfJ4zL
EyGAFcrYfT+9WTGAFU9zeTmHXryqMhUeM75Z6vtt6paXpy+e0HbniGxtnenLlQMGAieOoN84br2b
tmM4CLq77vufRkhNFm5yGqVbltXQNYQe+1QI1xSaSZ+xBypM34OjU1PRGp/Lw/kKUMTACkJ/L701
RfVe50OGWgVMoUpGAMnuIPASgtPcTgCIJXMGUwapz/EJVKDGrSjHNkXtF7X5KyJh/M1X9Y0s/0Fw
llpDu8+Lfc9eUGj91o5FaA7d7lA8goYCSCCKZ+I/5ovyLvsF9iQo7g1D4uizAoZ3YZNZtd82JRwV
2rUh1T8taRk76yveb3vCpwws4jEfKXRNwA9xnDaeDsB+ZkEuCS9ox3q+ENuWouh8fvbfyxyc3jea
G3AMKKU90jXjGnf7fIKVuNK+EwphZUo96kJFEVcQYU41Qs03LiKkVIr4apt00gZG5iy5qMCjONmS
xKDLeJnYR5YBRBg2ZbxRBfemI966n8jKDfnyx+z/NqOa+JN81wuufPClZLZkh5DRH7YmAenex5wE
ES/QFfdbBCn0l2vxPC+kL4wHnf/BLWgsJgU5C0Z07xpUq6A1LvLWLjji3f8X9C958pDJMno2kmPR
E+ZrwtUvAlEkK3DUy1NqLJWwDW4OrUgGDOo8AZT/DFq8ONJLW1+pHVmFv7A9jQDPFnQ1MhZlZvMQ
ZYYnUCSr86OHU5r2XtodK5+xj5qcYOgsFXWliHp77BupYyqNR/JwWvHyqKr2qIxOImFOXB/527bJ
tXO5IDavi8ctYRCyhyuk+hd3SzFrL2JB0qvBm/l2trVitH+JREDq0eNK0zBD/jbc5wlHQV7ggBBY
CDEvgVGgG04izHlc5IkC/6op12tBozAZTMjhYj+WkAQ3fOsDEXFpTNPVg5SQY6GMdQL41ROCPQQB
lPNPW4nravTpKpiv96BNCUSmAbJFeU6qMyfue3F5qf6/LwEt7/gNT5RGm3pHtvKJqSsJmZkIvHFV
pVri5HXn60PlF/9t63M2YVtsa7C2BbIrhFqMcp6fLfn9eB2UKST6ktzKoRnTjQRravTn+Ev+9Q6h
glFzgcZlvmqR2sNA86eBAx2YhbBWP3EhgyppYrKIrrmcYHzT7C88zCJyFvOYkBLJk2M5+l/wx5WZ
Wmw4ye1tY6m1ZbaySzZf8JbfqwS4qs0erNoYuxbxp6ggs3XSkwL1SoWDrWvIZzL0WXFFPvLhB0Zl
DW05FywRjXx5GnFVGfY2Dh8ZyPnKawftTzzd/HIi0K5+nX7QYYucxzRvA4BHx0oKzSVKpWNl7OHO
Ns5eL90fX45QAgATsLwLqLIB6AUbkJ7ziCaL/OjulJ8M2ZKKRpWQP2SIs1aoM9ZkMXO5XsWaeG5J
2FxSpz4cDOprc/fGMT/c/oecU1nx9WbCMOKDX/0FvljzfnYqGkjHGGXIOQkgov3mhgAiW8OgCU8a
bDD9aVRru01nkfYQyXqKmCtl8tdaG2kQBaeViTl+8tShOhyD3cCSZQybV2A/KIVQXLwVc5V7b0uC
ubIAOxIbRAyJyqQUx4Y8VPO/SqdHVdh10rwIluO1MJkYEIlrag2qb8hvSwLpLHw0YeFDVo1uMOVP
gFi2jkd/u933EvZLkNJpLq5ivmBH/E4qZK+Jmflz2dabyNPYXPqn53E5J7RfXFSb3rf9AdI2pBd6
N6geYUxnUvw7l/qBgphHn6xh4GaaZ0tDhz32YBVO1hbdJ1OoLX3aOGvxVCjdHlK1gl1D2McSQxQZ
sLhXBV0Sr+yygCwxpGOf/yhj7hhiuFa/0WDjCX9kKEF2c6q07MRpqNx3AnEMoATiOrKhDflaZppD
ibu2UcYWPcij7XPhwilWLflBUCSU6vxaFkgeXe7puV4rKj18C/aNGRN+2XgS2PldvF4LmaNIY4kx
S8V/zLlMhlSPxEBfGhJX4t7oFDL/3v1EMC/uSCkBZQX/noHRoXtE7INxbI/lJKFILAS3fHdx5M9P
JWTYSB4obYj1Q4mbtaLET/3hOrMAoF0QjirtOw3KbkuOS9gHsEZDubIY9LhCENKKC1oxUp6ipb1u
7yEc7fXA6T2KwOuhxC8fbY6kbvNJ7olP55niyFHiKDeQbDZTrtz7FhTV7z5457AndDcJ6BIq7yBk
VIygBS0GrNMN/yRLfxKzQaJNhtcn0wqP7RTkyhKB++MtpUWI5hdLdMSNiVRG7tHQVjks5xn413w/
1F7cYvntGYI/Ia3GFs75yibbNIuVz8d+o6A9O4oGruQ2/Afx34iXze/e0XMkvA09WB2qXfa40gqt
LDVO7GFKCYaUNkxRuyuQ4sjAAZrjTZn45lGFp3DZSPoaWq637Unqh3HnzX+5mbeSGTy3jmEiIu3i
UFkLbmwAweMPNjt8CN7GemBIVBxc9ax0aIDw0A47epEOoUfm/hLSo9b31olanTsf0Xxl5qXAOiM6
yqgyCBTMSeShTa3UpBWJojiQeQuiG8q41mrZOua83ZrdD6KtULSzu910KwjHy6fXZ6myW5XOvGGg
XxH3GYWfwDNhnD38LylmK/LcjoFz2cBk2M6tRpWtTZZor6ddfmKVic+QngD3zLp9djSPtoSG+jYt
LjHuLwcQ1e9owUmSUIy0sgPxTe6ABW1fhZdR0rx5bmhdaX+XJnuuj+zNE5iGVqvOqADwX3fZtUD1
A8qw5o5mv+Kgp2tR1OHNeRng6tUlUxeDX6uf2v/0hlm5jO9FgWNnKnYNL1Ggl04NI5TIFFB1Pxax
gm+vFldJSz9Fp59QUQmvh4jeMRWHe4tYBD3Kg9tNspy8wgXMUiaYcvLLv7vl661lUKVUHLyF+T3l
nivmAd77cBZr6qhViVTOTvyfa7SCQWbEIOyQJfo+sUuCeYpVJA/s+JDF0zuiA41WjrZVIYB6mlzU
kVgQ2ZaP2pFLAbG0QK1OgLwIUlWBkX5StiO1LVc2MH3CE64uTlQiixN1QJLcESRa8B9EXcgJ1Ucr
R2ipEqexCfEeeG4FFY0u6TMoiPXtRyIlnNWcph3sQgZ6Pr3VXjrDoMCnVvhrYUBsR2n1gHDEChYt
LnLLLMY0n6NAYRKtXuViip42NRvQsyL39JYN3A/B92dFIM7KuRRi3wRbFvqEQdJx39sfBbSnIp88
g/2vT+vxigBQd0R6UoeaWQjj10Jr8G1EBnpVDOwNWnJbBbwb98ZOeb2eIymjDzMnIozvVLai3v5p
CDqW74gpbYNsLUA1HcoVrc1LpBjbUJvS6ea5rY0/86dYv5v3KPkru48BNxv2TFv8DYU5BJoy5X59
Sz6NcRmAPJ0i7AfpmAhjYv/wyg3bF3BI6m/2AMROWUHXsIiiB+bnjr8Z2i9Z6i9tSDVHDMd+6Tw7
V6efrXdcndEKaWrfqj1L8WDtTH+oSLQxlorEAAPg12vSL4w+zeMCDrTu/FhoMjhDbPCZs+TXse8x
oEwh+6TJ0YqNEL4RtiYimYKh//mYgzgutVWmgjZsLq+U86jYfmKHUpMe9BBJnob7BcfuWjrS9s5b
5l4Wk0HTfNfY6GRv0UM4dCoasFYUJPRvXyXD6+2T5x3xZBEa2artJXFpfCxmgkFdYxWKqE7Mu1Dp
vzFAv8jhnzIOJJp1gYPVghPnEwhhqSvpbU/S08xPKNXAaoKSugYRMihSQQ10gQ76PlbB+2GGJUc8
J+qOgkoTnETo5EUTitN98KFK3yGXtMjuDymqn1QMiutMhDxm4Crz2Iq4j+0Bj8fTRzqrRPEQiHly
Nyp+YlYDcjuSNV/TT/MzG4rih6B1Cw9mbHUdzFb3SqpLyungIMnjP0y73eRhiKU+AqqVxPxls9dM
ojL8ueezfYpLOIZdvNou6L8UzwkMAv2Xxp2msFOB1xi/pUZhPCosJw4h93VkKCbZ4FU55/K0c3P/
+NnkoNns72xFyk6jp5DIc4AV/uwUWdp1Sm/uyg/D6EPzuR7KuAPV6HAoFdDr9uK8+InViWvkuXAJ
oV+1rFEt9srdVZU3xU8lliAF2AzZ7A4KQNNBoAokfrFxlLSTP943gPMdZO0YC8CpHF2tlq81qOH7
YfyeB2Dx+5Am/X0dFxTQVRl/rseSJOtNNF7UF+JTgbdXVx92Aid1vMVlunMpZBtKQIW/PJOYjuBy
Im+/L0R5JEF6mbuFsr2NfthDwpCwkQkjJOtksqLkxT5MPy1YG2BTlHKtzyrpxYZc67kPoCcvr+xf
342qlcYx7+akCafx4PryejELrRHewkjND1br9ndJOlmN0aPd1Y29g+b1ZblbMPJw84jLpiwY7FBm
+ZibBntqg1+FfeHGV/0iiAYPiHxlozV8Zs98hjRzd27IhcVCUAZQkvd/rabRL+dB5I3B/eKvaZq/
6QH/CRUDs3Rcl5r34bPntqG7nIKYjWsUsF+VrzY0ay8Wa+XU3pRZnOeg9/PuiJ7JdoYzu8zoc0DQ
mDaBZ4wdi1U8/r7zuMu8tfIClLVQ51XxZ1/ynTWFhzbwwqz3Ws3DMWL45TOOm+AV0Jh+UMAuRY6K
BLpDz1R2+c0L+mCRAwX9HB/Y/8VxEmu6sJd2NLFTX0xW0CE5t6zoauBFORdFCiZL6pnnJNEvO1ZA
tAWf4q4YWUKshFnuPMicwhhm5p2vsTTdHzQTfQHMTdXGkkRp9u9CGJc3eLJSJjl5+Yp1XlAa7Xr0
X9zG58DlCAqApw2iNS1DNkfM6JgMY/J7tKjM+DxyQuUBDIPR+a4uNDMNOJRQPLs4iwN09hWeFYDk
Zdv6u9IuZxTF0it9mc5GHB/l5R810e/42hchY3MGzgNiGSotBS+vLeUMklzYvqzc1usYjMkFWSOn
7PPXXxDBm0J/arc1dKx5dQ2klHBCWXDbD3WdgaocNn2h6UiXUXOymeIMgmELeuVSQZmzq1IZMZuM
1kT0QtSKxnmMdzCIs25BkOeRZwIblBgkQ8fudzN57nRNfFxTmEuoFO60RJZkLi55iW6joK6hNs85
WWqaTVZaSlNmcwzevqULks/wGOqfSDEyR8wjCdqNYJBcPBNdinwaqWOQLhy53gq34D6C1u/8mW7q
cIWNRteGvUp1qFrcJvVrykP13RXHtSBwQ7zUkItaRi1YM2wMK4+megJUlLPLzCEdU2iq8G+krLJE
4lQiYLvw/fUuKvHCX2QtALU+cwSciwhcJ4cBkLiTIQSM44hVe1D+kfv2f0/tv9Hbt07ax1YEbKib
3Yp+A4761rj3sC0P7wJLi47dwK5JAGy3fW0a/OdEGa+2cHiQuPo+lkwztmrKggn6UM0hn6uRWpC1
WFkPJkwEfUyHM1eJt28czFK3dpLLrMbj6ciuSg9EQWjgFgBPVkTtsxtWhu/U7yCiezdL9geWq/zF
hv2eT9rALyrazzPmjodapFr+LKJzLbJdKFiAn+KEyWsubjMuXaYkxHNNT/WlV8dP0AVYWMAzETNI
9XeWjNLXBdraGxOOf6RufopSeNqGNdxyVtcYUKfnaWWNewDhDuMqRVxiI+iztt3Gpir/GUC9C0WW
awrqpn3oqxW+WuXOucw1q8elUDxtYk9EW4QDL8XLhwEccs/67dqJ2YiTQ9Pv5OjcPTvZRnlKqVhk
J3jkTQHZKoGPwPa9AcK1zWqrqOESARibQXGi+zEvtuo+/vQUKzzEfLX4fUFwlqZZKpIKFZzPgYzV
EGQYGPMEhXP4EoYahddP6cqNR7N0Iei4iDIi5whTvQqrQteh7SvkjuZdryZTyjqfLr10IK/7QntH
eiwpjC7hIyj3xSYlRoVTVA/0EbROCLX58pppFC+2wrtBdmmrzJGyL9O7gqpkEtBY2SueMZ/eUBsL
J97cqhFoU0Hcvx6Ypq2Ig6J+uCJPeJ6s/v3kbujF+2IpRd989Byi7ryLFzkMQu52RPc3jfB6GDcp
NK7SX0yilIyS7S5R4wisWF4PCRSF5ohbKmsl662uBRqT1qL1DHNvdUu8Y/y1RVPWltnauWjtvFxa
UTBxZ5nZll17QYRBCNOK7sXn2vfW3Q7sPyC3TMcsyk9XekHBN5CUlkksL3fYipUHeK3VIwhEAFBX
HK2DA9juLccqj1EiHvrlpTEMW2bNJSvtVgL5+yKp/+xHJiJMLVmg+/PAZpIZz7oG2xwBjBM2BP2o
lyDPbSigPH9cDG3mR1TX5q8il8HRECFUDSjP47pjH09KZSd7QBH/Gw/6PbYk8C28S+xS1MnLHx6p
ZY44DIxAfC6TZLoB2K2ACluKCzXtFJgZcdB/KD3+Wd7ZwpAAia+d2zQILyqn0cZP7DywQ8cgqCo+
F3zh3r32+NebX4P8BVBEEu15SaEMt1QoRvKprEfK3OWU5/5dNbuGt3nG2isPQi4DD2TJ0qB+3I4v
mPljCDYFe1GScPAOXtYnMaUxNUNjOJK2WS88FBj4EhAzhOcsdfCruCcrcvBReiD7LmvRuuSJKIz4
qBYQMbxzDgG5ti6t69uzerhF+q1Huc+kKHM58r7KdSKhJIg5bZ7y5tlZUgDHtsfrTxMgRL/JbtYT
Ehv8tFj/wo7M9LqV/QH4z+Q26K+zZ6HHh2qKeuIyI6gZr9dfNGMcet4Pw3KLepasM3TnyowoWI+2
smpEZ5lOmEAuY1slHN4n/COqsNKvBhHXtOJoTf2VXAEzMV1MNOafDQLqRYKfqv7eMVU9KnmdcM+N
4Sy8de2L1B9QS+sI7PH2g9xs1cFsqzuSsJsyK+V/ule0SI0DJeSeAUwQaBJx81cl2essquDy3H3D
T/cARsISEHzwS/PdITwGEWIaGK/q7vLLKU8lIgpnXEQnvrjNhT4UjSLv3O8vEsjK6FGhNqsnSp5r
f1skNlNTS5HdQYtwi73absGGpKN2vhc+yz1+e8ndXAzqxSG7r2J6PzHe5t3AJIxAV4sZQlEltFCI
852ip1BlU7CaA+On+mW1TLcL5GQNCo/Bd58e0y7RFh65g2g46HO/Vo7YZGGHjxXGgeC5VXCunso0
BTuwPQx8JTmvwJQpfp7QvMsruWz+yRYO71YFRSk7YtEdnJhzg9yqpnEQ52UJ3a1p9zI2TrYE5GRJ
/pwnPE2NfJ4q4Jsif88xUHvFsuaJLG+uUmj2Hz/jxYUj9LrPKmQ58X0jCBzayt4GJN3dtRZl4G08
465Y97AbctxdcEqDQBzcYZscN6WW0rBNGgyEM82tRpuA/MdeqoHEqVIp3UHf8OjiTMigqjQTfXtV
zRwaFvy8vwtJpU+SwzCIojrE9OqPkh/2wUK7ewwu0MEQgwSgaduPSRcnOwkBWUzxQiDi+758f9DD
i2JRe+1MUEaFeYzNpUtm0LT0TizuWfjN2Ujq/pTftgQRcJVElbTP1r7HCuXPmCwYQtA9KsBqfwiO
kFnwmeIhVUjo/R/TWvGI1DmkKc3OqW45vx1izY1PESrr5JQTxcU0niBEbrLa4AaHkMHyTSXhvd3g
Ay0i8v5+RZJBv3DADwtTND5XRNKI1AKkyfCpqV52bEBjzVf7oOvT3U7XVSkJpMyx2jA8KquGMMAj
mEwgAthAlWmZwBm363hexr0rEEuS+msKAWtAdBVo1u83ynHGRAjBbFYFB2HihCeVHoOs9tfMnm9M
vt7yFb52G/o1INlHIJHcvNLUGhlH+M/Lu/noWrDG/OKrGi9dvtrWTnXi6cxRMk4fZ8efJBoSUuRa
/ouBw2y93rVMDkNm9rRqVuch6Yzpw7dBHOMsFGJ9cnvvtU+7LzKMQd7JuN7SjMjFoSa+q0jVZciT
Fx5uXiGLWh+sZ416dLHQfdJXYLTBTYNlA+zDDpZ6eb26I7Hzb0F3K2BSHsYSYQLwpoAhfHOBiyLO
H0pwSGfIuO0yZtoAnzS+Gy4rGMXZExh27E0EsqS2D6z4jSH+f2Mxlf1K3a/5XO9sx74DUxZnCkcY
7Lej2L1nv7hrDAwKYbYOwYOiJZMAE0KhZsh7x21Kbxj/4RJialVT+7bA5cWt5/TqxtyTObLhpte5
nF/GJoCBLOky8cQNUnH1ot62xh3GC+H/and4C+X5irGc6RXjqHXEqHFqo2ki155WkQUnso1jlpZ3
UBcxi46u+l0ZDfLuk/Q8peF5nRUY0pYhEFupTk96Ydw2udouW8b5xb1wcKBastfgfz+0YNef6uRK
a5GLgzEeTE3RVz2hlHk/+Xl/xWevddNnXKjO8FJPd8mzVR4uRYvLntFAK8RxSwm5NsN56J6UhaRR
uWHpV27xGb8o+gu9D6Yb2F30icIUmT/uAIyeHtsXrHNkkh/rfIsovBE/uelU95DMIn8v5SYh768z
2FVB/J72gzqcQALOripJA/d+QqLLVzvVVaSBOFO8XGBxSSoirlg5lNcltEJDwIQn2N3G75HtsesM
CQi5/CB3z6EZFRt76QTZl3WRYJmudQpRcuA56EdQkWNhi96BooptQowZnWQ/u7SkQzfx5hXpaywc
JzMcH0txHQhYXq5o+5x6TMBOq6IVqqZxMZM5uCsoGruu6IN+1FICE25e2iBPhDRThBLnDMCR3fTx
hyKcrUWX5VKBHEkNsmk1KnKMx5jG5Z2h4389aKVz13W9BM1rOQN8S2KO79G5qCX6coszzleHOP4L
E2lK1xfSAJAHkVJR/yZFhRRMsmgGY/rk1Psm5+Hrh7hPoz9oFd3Rc786B0eIEmfIONI9zUSJ/dwp
K8JxXw5CivqLEQX/GZags6chKV8kkEr1c5hzqqgkMUaaX+lqQbJV+5qTwDP2PFcjLZAAwUEYbzuy
IveuNMEodUeqfS3MUswGbx043i/4sOCKnk+JLL5FP90mrHOohcbHnDnkXtj4H0m5dX4ODVXLAZZ/
tW7yZqEcLARbFnE4e+cXzPnd2DV3hHjXFs3vQMtY1p/wXy2q8+C1U0Qr73/uAZx+M3xxIwFTCGH0
W3BvSUh7wOfV+EeCzkybbe5NUHfsp2iexfxcgmpbl6Yf95xOUtYM6buI3Kgi6YOybNMtZNsqYOxh
TrZ0p/vszHng8hV4MKkttI6U+jpuDFljq7iZCrub8J0bVREHRlaamYBpuX3UdCLGsZt7c0sBgsJe
F6iL4+GX7wt/RS6kT0Dj8AMPGdk2Jza2Qof8bXGz5TLWiEfSYRaxnXAmeOcBuN+WzSIvbR7W8V0a
BjAteylDeoWyq5W36xfDXkJsxOh/EWKvcHEUR09OITpGNDt7pL/WlXLGjaEcr0aaOxi+h63ynAtL
QG6hvLFqpL2vFq40en5eXJIPzIe5YvRcgWztGvDQIrwFWq+KLhGlZCKG19NqB0aDMe8F/6TlsE44
qRKHw4FXFCMjR/6NwzZ3yD2OblON60fhmyuPieN50R1azj6G48f1r78WyKTghBcLlT+gUkgBrBuQ
CSKImqZ7q0tgz52YaBVnmYNQ+AIi/hSoEZJIgj+biYbr/Y0hVK/A7NQCcCo5w2lBJtolhc8q05NU
9/dXh6cBA9mskjugDaz3Pe5yQPq5ui7ElOLhrfYOs5wk7TkW6RS3lOIXjaLVHfZhYQgReTp92W+J
HWhPIkxU6Wgs1yr14bdTSqg1kdEz8vL2EXxQTyB4kaTlbfG9f6u1BsBCsMJjSNkfMaOX53DGUhH+
W+TbkM4GV9FZnA6xgOZJhJzdB8mj+m6lohZO4j44yv7Q1S6Oph/e2Yrh7NQr9bJTnEPdxPRU2LNq
jzp4DFZy+Gd9oMam51hOF3ouGW0Z9gkUVxMxRbsgUgjovKYpj+x0FvKfmyUFEgQ/1ZQ+XhGt65/e
/lqBOORjPlTEcVuN8I1uXLS/gTDcA+2vOOe3qi+IjT4rwyM1nSPYmDYZPiW8rzH6lkpBwpkyECec
n94EH6S1AEI+zPipZq/WZ90+A6uGtSGthhirk9bzfxXB03qS/uFUEF0UwughzRi0T2JhT4eQoz7/
0Jlr7xs0AEBrZfZWCszWi8cyMJU4v91lyTwD0XlOhLG679fdTFAJV+KSoIUe1bqMP0ILnfGI0u6N
m2aD6UD/mB/l1bMv+GHtM8shNtioxaWU7vajiygqX+e/3nxajwOx5mq6ffbuQySoOKsxeTiscx3p
K4NA8TvIIF1UylCcUrn0KogHWLgy/Sg/TLfInDAmOGbd2urHxC5UNEt9lXNOuHKQR2SqOntArDAI
u0xR5sqkbgQHaFpZwmN74QqXGk8By8JxTnaf+27ZKUblXEGjGVCDEdSH2KhdQ8XiUcDLXK7gI5w/
x9FzdHnldei2+B8O73C/QRhWdCsXP9u4F+R1HLohqpVX0yUzR3WnK4jXiFvOl/FQVDStP3GDdlrR
6uy1Waclp42l3kN3pI6bJ6WEUNAXNAXhwC7AGrLVcQRzLYm6dbtnOr61QOQTQAlr/SN+HFa6ywE3
QOSBD3Ht8BI9NWrvfDYJH0nS9x3EtfYw5lr9Dxx9fviefq8gL+xbSuyOsCcIJOir2qQdoXsdqyqO
0hkgVM05gU1B5wAsXNMepDEBF0l185OpPxofW8cO+/iuqaskoQOjYdv5BeTlGqgi9sHxln3KOdX1
TEyFWqvVcb6x5c2+moOCYbiW2RbbyNm6sLmzMIneluTbNJrR9YyBUkaCRG+gblM/AJHZ18P0/0bV
4O+dIe6HacT8rDCqleTA88R0tXWPghSxH1ibjPM81V2uAKntw/zkSLgr2j3XXTFceQ9ssjn0lC+J
t+cZElSFMQ6iwPstemOOal+tishweZIMpuRfxp/vhhnQVZh2sBHfF3EGDMfVHqIwfprISO+iaPUF
E9QZIAwU6ZZykwZvgxo/SY9U8ZZESmCM8VPamuGqobQf47uVENjLm/tnUu8t/OOzPzAz/03Z4t1O
f2oMWBv5frafJTFQbU9d4NT4c168kOTfkENYbyHhIjgFRIg8ednPdVGLVdIeTrEqJifa/GQemAUk
3gNoxWGPlR+tTGegLBkxmUoyhnHK372xEcwSDKZME4oYYEDoHM0m0jUaZYguEYCY5qmR5p2VYAOZ
+nfoupHa0VuviKJN2zFpkNrydzdAmXzSACXehqVoPF6/RnfF3gChB13w7UvRtPNMbyq6V+zeyjYo
yU++u+Zp6v5g1q76PIZ2KxX+aIY8z+fOHWa0NnjoM+y3Ti+A2XPlFGVLVwn3R2VvpIwuPOvP4ddX
WITS7CVgmjBWR4Q8GVVaBUJu1TrAFvOfq14XT+Yimnir6p80Otghm+Mg30vs6pdZzJXnfTbGY1No
72GEJakiHl/mp2oB6KmED8rc60k1SHrxlQtsIQ4oSN8N5CUmOD6YERtBUqz4spJK1VAu1PsaHpT9
K0KpHf+eDEs/LIHjQb9ouICkpICb/PCNLc96B8pPEIfUMKpRGb9AQmDRm/r1BvfUIeobwTmWKatv
bOPijAr7Hyq4HDaYabwWsd1KKDK37KtRl3HxfpT4FIHE0+12td4Jya47DDciBt5ihAYAvOgm4k5K
W0caXiyFjz9DfOWFFcP4g8GPBVzXyiWBVdyEjhVSj8s4YXtjnS5QlTKSeaU7DCIUOy9dcivDUgM3
1hifH013+00DPRHQ4OzxwZVoNQpLbsPzFV4IdeAdROew9IZQEMybfrZJaByCx5SrL6U/Xl54IYaT
Fn2T1Tp9I8qaeE+XAmI9OSjt6uMtrHlDztoS2tXL+DRTHhXKGFadzQcGjvcDXBEIuHcDgcWdAvf9
AGrXYj9l3yw+fqtZOe8sS5rUiPIslp31JMaEOtCYBzziWzGZK4rwzEo8uDCtS9783XVLNVHIZCdn
nZ6qSEeCUrBaiTSMrXAb234ZqQKBPHmn6uGsuI2xBY8Z1oyFK5zK7yWkoHLuZQzoozFiKq9epHq0
WntYathJDs2uz7ZIuFKzGRtp9D79TtULZUb+/SBRlN87q9JJbF9z+Fz1QAyJv2fuTvNt3h29OV+U
hmpKLkFLxXEENh21IRslPZh8krTLWQNpVkKbNvNrSnhtwXBjjusu/Pb093vQm8Sp4RRzECyFfnoB
Y7tGFPMG55klQdF6PxwfusPb+FxBKa010xJ3081lEBUe8r04g/OAtUc8i/ZRDSH9nxwUCU7pP2to
3dUV7D3HlOQeiuGFXngD0BIuwqaGrSgO26m+mf7K91gzsLcP7+j4HG6uJW59cIMPGr8/mCjKE3c+
gQ9/+ZFqke39CSrI1uG9c749rwsqx4r1BYa2fVjpbANUSwYrrHgfKF+fPvuZGm1OmuOjJ4DToMBG
9Dz50t1qZOHdXr3vuLc2BONQWXaml1GHjGc8Cxf0gECPCvhPMWAqSWIN7aer12kI5mzoZVLemMXU
3jA+9HA6ttEi/UmGFS13HpiBqpx1bwUHQUCHNcbywL6mtsk+XccseH4OgWbs51vXL3Wx69N946jk
k/9NlZSX4DIueyndKwJSigq7veshSU3fg7z9R7AnOCFr6ekflvlzhJx6bG/5YYTYKFaMHR2dGnPy
KQx5d0t40DPb8W77SvTNlTrvA8WP7IZj1fT12tfErkElUx/dkr2h74p7T72p6K/fRin7eAXSgE7l
BSJuBm3tocGITy3NlAUwlR3o+y5TC1iH5xZb8IcZUmNGYVHKY42xMFmU/Uc5CNESIAar+oUmY72h
0mUJrIT5oD+UWisvykn8SNp//BmyS/fGh1TdCVmK86QjvMNTE2Mh3BFT+O+8sc0lvHKVqrd4b0R0
LNiYG4sL/BdGOr+dMXo0c/zURJ7z0KnwA9i9ShvJDK9UgV9R+2u8aKj3gVAu7WTOHuEKW+kJKc9H
ywPIi2rqZK+7/5uoWHgqFYNNZfzebOHicx94cNlnxN97tbkrRMdZa4/6uyrnnh/BmQigQKc+WdL2
+qCVOzPmitJ6qToG/9lRCDZ7igCwc9JUlQoRYJQ8+zTZQiT/QEjfc7oXfJwoBn+Z3PYPPngMHsLN
08nDndkzScnNeWJ+Q73uqm6z/GUBiuIodsw8dPNSwa3mcYnKblty4WdQx4Ppbmamikj8TKFcb6X5
YNdoVbhn6SwEdy8ltM4Bs2FxjARMxyqfUrjw6xp9lPpiFxpPx7A0j/KDgl5qSb2t4IOOOoECVJfy
u1KZbuKRit5fjPIwXotuemv0Pq5AprriBAqn9q9+Rr7M03kOdU8RQ1TAqAo1n5is6bwVMJ20auhG
37kCs8ULdEV2z3hbDblQm3/BxCv+a/nziIUXSRSrdzoo0jjlOyGeqgkYyL2o38tnD0rdibdphaGa
mTwbgYzY4TZ8mEOBm8NlImS8SUF4lcCWMuh1uQtvMbOoeDQtpRR3hWyycAzHX5wbDWG7btExXOdw
sOTntn7Ozx+ts5WFNklT2Tw/RyZYex3j9xZmQUaVSSKYczoZIFNCr9MDTQCz47Tm82w/rxWhzv2l
g7bk1WCIZ0IhGGvb181C9qiz/H8d3TgWV35O3uNaGqNVjcPN8M7claBVI7yRbctpuIvl51z+n4mM
vYE4UfkYV2BwNmyzgmSlskXH20NAS/Tgg66xwcJjKZ2u2lT2aaQD8ZcFFg7GLVHXi5jQzVvgKlOw
c3avGVpgX2KonxbsTpzgo3/icfwye0QbR1389ZWIifNsFE8By7OqhcR7n9pQDL3PnO3s6bJIhbfI
G+rP9jKbgWvpYYjtRKUpFpado72fZYJNX01lDGSSeuCW7hvbEtbaSCZFf53UyalL0cTvez4awxTm
OF36hT+slYuigv6ajiUcIyT6sCzFvq9p/wDHZucA0dg9yYCYYEJG06AxwiqKLMvLLUZ/Nf+FSlRZ
fm5of0d09fED3jKoMdZDrOJSqlIan7pzfjB590ohWS2mzRuUJta54+gvf4/v3HzHEM4WpbXQrNeT
4B1sdon+ue907+9ol6229vZpbnRy6NpPXW5Z8Ucju2Z/pmYYDwgWSmzsZRmUPV2ybA7ZUOf+Vrsj
1AAWyXp2UhFMzGhEMDw8hGExgxs5OYJVe3tzGLuAG1UG3yhrnLQRwrnLU9o1kPYQqiueUlwHpMwI
/2qw2+sE4alIrg/+dEzkLKDLsf4kBbkwCv6KzYI0UGz2ZQfjf3CHtkA7+4NwSPza7NbDFuK5fJS4
XVBeQrtHPOQBqHbLOvUf/db9cUtxYrpUgsn/BsjwrzfIua1vlnOeEvwrDuXNmyyoiA3ryTPNprUE
zmU8F7ITokF/iMSBaxE3Dq8Ew/TtRh+L1hadq7QLgWPDymVlEpG1PDxRGe3xzPS1WEh8mWCKAI8X
2oK0ktAuiQhQ0e1KhkVIiSjnASndEN7qpz3jI8Nb4bzkw6Pprfwp5H7ckM2ksvgIKHKecsD0cK25
3TbRbSD4Bu5a79BAR3g5peiI9ARpgvDxvmTdMTgkk83GDyvzN4XfHWU5aNAH0L8wA0bB+um+TP4W
unN+gaTMas910km8iuVVx1Q//YVaoe1p8zFr5uw0cOZ8oArvhpgSKdRxJGI9Cj+fFogXe1bF/ZFg
hKj/3MiIThC62/3fuf5S705DtRn3DiImUasTMhJWR+lSsZf87QB9o3j+5maUDFlMMxoLV6YHyxF0
UGBL1pD9RQrkxfvcqUtxBmJE4cqA2vXNHgKufqKcpu3XokO7i5JmOQgtQm8OvykLUp3PKHx7G+Y8
6I1PtE+Ca+pv5nRHyyWYHo1Ugy1zrXa+DoRPW4me77je/7Am8AHCJKtf+6nj+VgbwBFMYtFNw4yh
pEQjMXhqCRaua1u4veL9Hqyv/adE4Ncnv+W7Jhk84Hnq3n7w6ciHj7QyhcXpj6MI+DxPuq9Uz6h4
2E7fCJiCIXmR+Yw/mtHJhML3xUv0i+HYxsGAR/ifWIaLnpf7Ij5Ane6DqtYq1srBw0blrk8VyHUA
KXU20J+y325uEX4jQf0TmatXqkovrfqMSVzpbz635gv9oGwzFTVlb7YYyjveVTczMyYqRegHC3nc
ONQMd8kYxtQqNpqLcNOJUuZmeZ6M/Ufj17rmwHrTDp8Qv5lc6bo9InEDu975PI2kTlSpU4nDiXBq
Tnd8x76dBEk/HBeHr4napQbHpkVufCBJqyh6SFSHdyie5pa5vZOMP6NI4NGQ/bsG7Grs0iTxsbNB
CPRftXYP+xqb3tWjD6uSzngnoaMfnpdTGxD2qM8awPGmQ1DyVhZo+95eloAv8f1vlvxhcWwgiuYI
w6ijPHwF1cJ6xMJQPjaEE6EFPtq8JZFq2YzVw7P7dvvIy5wtypnVXK1uHUyG/Cb30IcYNtUXsY47
hhDeCr+MjD11+Gvw5xvYRPasIBDLVDy7m8E07ijzYTbHLxBUKD301JFMPezG/UJnWJAuYbijDNFg
2NXjDXtB35WE5JtsRc4v9xnmoK37N/b5aDyFFpxCuE2QOrpmgmMvydZTCtomxPK/L7V2mMW0iCRx
Kz2uwbMoJd1IWWWsrN5v2jQSNvsqxKiiDi7yd2WXy70HHRMNpi7TTsVOnaV8yJFei7Xp6hdyElhY
d2ggdTMwQIjTtnb5wHKpKs75kCVIBpCXbJHXk05/ZPFyZ6WBp+SrzPTPeO4/dxgQSG0bv7fxXFa1
IBCcq2rjETv4drKdqi48qxRo4WzHRehdv1rlu5lDxviAJBWuvOgtiU00oRdU8txjMYoksvVQVbMJ
3LCbAJBgyksmLS+BMfpdS73tsfbN4w81pQV9nJnzgwWPdBkHqV/LGLIvVKIZ9lhqgFWq40tUh5c8
/MOsbH16dDyODWBxJ18nsD5+jTcnhZFLVBPObw7y0phQAagxYcOIzvjmNBcMqQFynpI3yBFN+8RH
LHNLZ6jenNAscNyCEqi2wIamR11v2Kd7i3i6yTtTAZmsQKjdp/QKiY/UZtbxXDp52Xq70dMvvZCS
RoQZUEuqhWrIOswUcNZd8j8RoGLQCwqfIWlfeby3cFDS7UiVzywSSEUR2+unasahR13unLpVfOVu
MMpaSXqHJ832BPvm+JKBziv8O4qLKejXryMugVOaUVFRTUQhV1PkYtHiZoXLKRM8OWK6T6zzQJFC
pq+v3Lwo0Za+sFy0BfJ2Bh9QPyYpdH/TtJGGTMkZdlhDBs0rHZzcumho/D3/wzDstO8ZfpZslKo7
2MuewkeAYfCkxoCKqPZyKTOEVcQzQ19gX00asqw7nFzRf1QMLVASYGONBb6+iPIu24zfcbntz4Ys
0oDALF0Yqc+TyL/e/hEm0I4dACLnXDDgadpUdBteSCZS2VpVfq5k/wmUbjut2PGSXQd9DAfwYr66
khAqtIo63+/TSQ3D9pTLS5Syyos9QpGLQBRt5sGfzr0azYv6+i922At1QLi8BPxkxTGdbojk+kta
PHfCCzmEOztnCP3dZZ6ldhoV2e6hF1KQ+jZmjsfE+Mbl8ULjxfKNVhG4d+JuqhsGQ89epFksHA4e
g7eWldrkAbRRfaVnSZsrWc9e/OZwRI15AkoxRQDnp4nsktnRDEUob5SLiSLsb0eRIW+cZZ/UwL2Q
312WiJCpVgOhqxW/1cBP3mKqsR2qS5/Mk9mX1DPEq2BzsaKIQs5DBqImlSLnPhSDX9YTRs2fra9v
MOluG21ov/gauJZ3/FVyFr+96BfihbE1T/jvyI7tHof957tJuIdAudsebr84UphOsXkXErhLJ0fw
TIrUO/GDMo3j2vtwD7K0X0ZM/y3o4Ckqp5S51O1BU/ur+llGtNyVDvuFtYPGX0HR/xzdt8QHXXcf
/g+jtWbLLIN2TwRC8twKA3S3dCwk9lYVvsdB2U6x0Eb0rIXC6oOtHnSLs10FdASybudnCtX7jKsn
K3U09CGtQv2C4nluQlCsBjr0I+OjaicTCLWwxTN1inTjTUL8kpHi0DhRRwwVsyHkYAz9zYSkivXf
nboKUGzDNTT0RDpqFpf0mNJ5/uTborhau9K2oXvGDVipSozXPnIHMcUxIA+JxlGayOj09mC8TEqJ
7NbeOtQVxN3ffeNmyZOMRVOCQZlwXexl+imZ8iEYQY2reuOgud0h/xw17NZMtljh4A4B3K1OoDKm
3YatGpdprwZWA+nerdlWuaGe3wwk3Xr/WxSRg9ZnisiS/ZKnZtEV83tySz0aNxseMDrAV7o6Ipbb
NX2wRs71PWMgoHOWtEcuOgB4sbr4RF4Nyca0A5ckan8lbAoo5MrpmAUQBa1OsYOedPmoCib71if2
/P4MgYaCEDqr7UmAJv/jXE3p273Upsp6vdOYOTTbta6gvpfHb63TFP6ZEGQuo4Y0Wl5hkB/u/bG+
y9hZPFticJG6zDZttOJAXxZh04cu2N6GscVy+uZOI3TBV8ab55hKiQ8CKjQkJDL+QmHjopfcCsp+
nqpTtBNYQZq49pCzwMj/G6Wz4y06CyZpITmyzvpdxkpW9cO/oH/oKtUaOxbB/Cq5KaIFhmPDO3q+
itmjoPN9EpSBp3NvNohRFReAp3K7OdGwlUuCn49NKMQ5NCXp/d3eoeXucfxDPXcmBRY9mUCBOsH1
3GIETbA0onu5gvBOS9/8Blqa/gpjPKrsYMtXbqFaqIZOlHol1jecWhxvVNB1ygpgRbYtLvz6mNFg
A2LsborLD0CnHYUyfdO0FYasUBqBr9wOomKmx8h0OzkH/3dQo0Fu4VDArDGaQt8f/egJpa/+nwg9
rO6SSQ7DUtJWX9LODnylR4L4VVErFZUokFSlnDL4qC2HbqDoNBA6y8Mt6XMUooPnz5nkKtIe502C
dsXS4+2KB71FqyFZi34xqeTBxuvaIm22wgoVRzkLFkrtLud6/sckHhOODBn/3SyIjW3PttWSRxPW
4S747n34lxsKSsPk7StTmXdy3B2zedYeqSul83sxj05gim5CsM7p/LzA+wg7tGprDhHjrJuHjsWL
YZuZnDMC2lJ4tquz4R9nGbs8iW17W0pxUOM23yoDI3LRDvS2iIlOLmB9fv3xXkLbRPl/hO+cn66p
p5+ZLp6FLPS5HG+Fv5mpBNR6SV4VqgSqBrJyjecM9793z5QfAWJ04j7DYJJjq1Bd5dbVGDXOtuEJ
9KFrF27l8wrm9LNIZhj1mq5UNxTRZEJbwFTnqbxK1Djr3SWnv8FZvovjZAfgDH/CGiso9bngeria
W3NpOLgk2iN+w8T7VRUkuOdoDMwAAZXue3plvdRG7AiT2zWfvhcE5NhmmH69cK3A5KIfZ8tMHBnI
v1vSNqlvxOAOODyeLY3jPA2gw5jMBYBEFUGEVHREs24w7jG50dVnRSz/8dr+s3rnVaQ9XFmjRFxA
fG3cA5Qvzrq+2Xee1nl85kwzw7p8wAEtEmZkRppDFMGwiHV/A5q09fUaIRXo01aWO4ICevCql2XN
PYThieeBluDEq5eS/ue6Gtid49IK7Snfnr0XW9A9Gbu0Ya8t9K4RN7+ZRgazQ5yublCh5ENRssOF
xzuqCV28kNzW0pfwuUCsDeGmU7aEgwxW0n4hkQvsznjIXOfWdBd8qYKPNCJgSHLh63fEOVDMc84d
4pjadxtcA3mnK4iW/4A/BkRRfmg+ekc8sEuJ/7o2jQ7f5VXPsGLHcSBTslgOtBmz3DbCftH8xv1w
XTaCS6XWK9tgT0OaQFA5DGBvwMHkii8YLQhf0MGG8cUBp5MlUVcG+DQ2m6IyDWmWg+ajatmTC9Z9
MZcGnJ14gnzPqzlvJ6QnXH8jT7UKQgfF9kayt8dLqzmaRZ6COnGhx6COHwn5l8irJso5ty8u5Hfi
EuxBluJc2A8U/YFqaIAPjUE6xPtKTwLPieLvk2T8otH3LNXnpMFlpRpmJTEFjn2dPbnDFcXEGJdo
zJMn3rwyadnWmuSHyrVMeJ7yLmcF5IbH2MYpIeHXUlFBhGPOegNB55WgxSChibjxGTHId8U3llct
wMLOD0X6E1AkkNaaduIWo4tN9VXevsFD/t2/TFTBzjrtN5432QthcvSjOP/RCs4CNjDaOeMvd8D+
Ac+hQiIbGj0k3+O/yLrh4BgOStnG9cjdcBubrotQy0RHK7AUxIMybBLQSvZZdjwblUWS1QJ/O4qJ
5PpQsH1GiX9DNazdaWYRQhMKjmVK/piYf5S4iRKvNO8orBBn7ieVdK5YxrpUS6Irbp5n9sPXocf4
EOUulXXn39oULMVhfs0cfynp3Q61K9aynw4UAsyvLibUyIhn4ixZhiIdE5Ph8Q9+w1rcsIoPik2w
s3pyvCK1kFH4qcj3447+zwb9kA8r4dw6TpTzNcy/xj1au32PfYGGsIvD26uifUdsx8WwD2gjjE+4
GmMTLJXbWFQM4KdoGQSXdd/Pt6HeBLtPMCJa6UMoR3u6fy8Pch8S9AZKVjwgWOY7YnxmoV/1ZZdw
2pUtUw0jJXHafkPtP+NYqIzgslvIwpEnVz4oQLkN1vgt1jRDCXLD/ml89Mr83kvFhD0atb1Tu7JT
/Il792nQGDBSyzcQP9USfHIKI1l7nBqRiqdQLhFARur+OZdIsOdBiG/YWJil7MkhCQxMLprIvn9F
EXx+yBYf2UzqXojIUk4CF/D3rivd4mcjHxpSunfY3ZDb6ufswnDXXaIhVorbD0orezS+vNP2rs+y
Pt6Jxs3I80Luz5xzA7AKoiCs/MWu5U8gos8QwOXtb7WT8bc1KTmk41QXNpFIX/S7PW+drsgIxK5v
bxauHkZmeMUVXDBdsQYlmUjmI4TzeGIujC2s5o49nnxXMkmmQg3dPXurQMY4kvXuVc8FacZI0+yI
OoU3dRn2dEK7VdF1d4J8RO/kimpLRTdNXNhecgvO6V1bLrkXG34gow7DthypXQK9Bn4vp/rtVPk8
F9A0zGOik07f7I7WjSswCV/naa/F9y44nRzvXZweO8iPz/HvZZP8lTL7uzUA4l0OEvJGQixw/Mku
d0wW5dYi+ia2/vAofypPfNNoBsU9edFM2m9SzeqzFPrII2nOAtdiRTeLKLipwdKKddOH/U1Zv/92
aBURHywLhUH5EViBd0BObLPeq6yPxM5yuFmsVreSOAO/xxqbeOLxPm6UILcdKxd94bHaZX67kPv+
389hVayiD2SrJsu4dKQl7bpnsk1qn41L29wBEnr/d6uo3zAREBpdAgEXJtjphAXAzQp/6TPoOVmg
q7E+kdOm+Nq/yLefzf9GdETzbfQ9Js7NAnBIvzuAOVdjZuZuGgaWnyHuz1O0UwWOloBMm/ihSnHO
YbrjShLFxrm5eg4cDNOxYZZSBv3BXUbHjQ8y+keszfq+uSla4urx+nNdRw5CFzIMTNSjbJMEQtZz
Z+4LgOi2JvJNpdOvXWxclqQy3bHcEb0ub0Q+fUTQkb47hFUO+yaI5AA8kQl+MUydnIJcrtkYqo0r
hhQv9Q6FhptSWSj3u/Mqq7astSJocYNZV1oB7hgJSuGauDI2IB5eoV5DmB+v3z4rIp2ldlimsgSk
Uu7NdwOmCd3ZuZqV+N2UAfSJhRSNIiJk3XpeaBWpfni23rsx6FN4vhNUshhacX726cenVtQU5p76
P8+QkAYQahbIJ42LKQogM7YD58NoOg0efPb43X07WqbalxcotcIsBkhO+lCRILp+zV8Hg1Uv8wTS
hqfEYmR18ULEV0OtUwKR7TfI0w3nsAummB33KwP7qXblAi9SzoA07gO+yjWAAuNsssb1PfL7NYlQ
SAJzaKm+gfLK4NFcKi6Rmv8skK3JL+l0aumNnsjWjeMuMJuFsvPgYVg6y90YpEFBguUyrLmUahzn
vBngg8PDzRHtvwfwf+OZJA567e/UH0CDPmw/QsdGXT/6Dj5szdJYEUpczb1cCrG1Hnk98rUq9AxJ
a/VtCl2hOKGdb0bgAvlgirBrcMzuylGevLjO31GozReCEUPiV1bXrm3DF0Aq5FXxc6Mju6bUfLsI
Mq7McxOxLPTk0VYZWThhaD4/TeSxhSEOaEHQup98JR25jrzma5qLqXTnaqdxnVMxtA6ITbP/EcjK
lgKVoRjDtDOjQWNBsaRPmT8i/lBWXo3lguWtNkNGh0Nz9z2sxgFoqy23X3i3rtOu72A/4Bynncen
zLLCZ1ZN38fJAmaTZzvxrxcT7PwoXW5wmfg4ljKgePD6yNXL0qHrrqja2u7zEmKfkmH/keKo14Ux
OkE91hnpQDAXw+qqh5aiAKQr3XJuXJyVr4BfZX6XqWp1+kjifHrGTBvHqhTK35TIzHT4xDUI2KUK
l0laco8xSKq2JXXgTJfjaVDMtLG7PWhHK4IDXns3i0bvPvz2HAsVbXgGnKyC03u0y1QAeroitYkm
+PCkKFS9pRB3hU5RXFbeo3yYm1wpLmlWN7tGiDZqd8a0xUbNp58GuAyhZwh+/ogX60xsfHI+W6hn
xhXRKpaykmaOsotDPYl93Yar1fEEOZXs+FZpZhOaz8XQ1iv8OStZZxlcG1GF4U2gyQJqvHM6ZfY9
8D1pFfAcmjVShwC1kJhKaeWV3fzLr9VZWBwdO6o1VAaz5RRiDNjnR7Aff4ttFKxDS2dVvwamgpOH
M2S7NF/TZsBQDiVKNHZRCF8sx/02RGvuAbYoXzluqTJX/u3jRMZXp/EfUM/8wyb3MjJ/Yqp1Ikmo
Y9Y9/j92VnUmFYEAWLYMAI4RQ5vGUvZo2ktCZn4j9WWVmxEGBCNujyXjWddoT/Lg8ncj5yHyTssP
3GE1fXdNinj/DQbTKbSfrdlB5nnyjfeQP3olkrhA+vN4eGR4BfB5CoNL1f2bObzaj/uDDKmYHKjp
8J22LeeNXK4bwoWbqzFc3S4GELGyfx+bSfIwu3K6X3pvhtg9XQiy47WmUDRywfbHZzSCNvzDKESX
7gGPhJ+n+EJfXt4aExeY6PiqPDKV8mPaJE2Sqt+HNw5wCRkq1GWAMWniY64OS4jr/Tg0VFYb0bTk
cH0/TCySn4nqCT6bNZ1gm112dBgMLZYhlRZhheUblaiV+RimCFkwQ1dbDWTpuYPeU07Oui7eGd4d
wXRkLPZ6NVvRLoO/vPHb4GD7o1AYUdZ2WD5SEk3t8Jaby6hEZ0RcUWP/usB0xRsS5rkeEoOsc2hK
Lnwv5xbN8OyGIsm7AXPmBPaUB2tCKkUUDbcPFCnmumex3G5W3hHTw2YCATB6X8YAloMmote/t7S+
qp3JiR/ThkoobuGOnaY4AsMJhtfBl9ZKtyryUooWDLaa2r1J+O3MpmBpXO20ALr9rLdgluFgZsth
9jzdlOitqkLY+h6Qzk7Z1MuleDQUoZUsbyjSL7aXmsKlYvxb9NSXg0GkwHwtTh8n62PIiRZ/0RJ0
lrDU/TfaQ/VVdghR7DPq6At1eTDScnDGeGJLZ3Gigsy1Y2sO3ixSBLIVC1LDmWWpo1vcn2ncuWU3
7RpCt9RozE2QI86/ei3FSq14uuJi71NMnWYJtI5f48nsx269ESgBu9zOF9dm1SmAYcHekO2TYPwH
LJ113S0vxWELmJJ84Zvb5DQigBF25zrqzcKQiRbq2fwi7a97Q6qyrpt17HvTMNnDmRTjyKH17ylf
4B9mWQXMtf4a5OQyUYG4zKathccw3C41egiKZq+7oNRPoZKOCO5B87sA+FyLYZf8pqrqZc5cjhPQ
Tine6EX+MAyk2LPbOPUwP889zzVzYQ6sg9gDvDUts9jnQo70PpUX0QSkSGJRLifdK4KCYC6v2x2a
+bvpEauT34c7j9ofdvN+9iGjCxWKta6XwbgEXZh3RFSyeVp1Mu3KzU+Iq4tXXHxlylhZsVDuKjQ9
2hA2d3XjkoxnaS1oYhagUcZfzDNo4+0HHoBvvskRSnANmOzngagTFSbs+sFG0+mYOPu6GsIVhQLY
DSEo1SsDa49fsz0yIojDHEBSgvRgfxPJUIWGyJlcoKS5+oDisS9bK3+HqOG12F0FQQx+/GJRuBB9
igxZAP48epxQ0Eo6YcAhVhihJidIBunvFIA0h0yLEpXPoYxXovAUbUlIHXB5cXBeJEEFV26LWlw4
BRPbG1a1VSyLvLLTdSemy2DnyEUKxBJir0FB4LgBfKwRlGrbY7BKwHWyRsBhzp71yt9WCQdrwwpE
lgxqeM72ds+dftXR2IkmijDBgDx+YPsDF0adEGwt9wRC7Q+dDF1EEV2BvtTSNSl84LxNQF2mKYOB
+CkR3VVGFPjJzRaQHyvLv4aWbYxTJbQnalEFmBeFjzRjIJQbYihZnXBRVNIyVuEwLVXmvVxEoz4p
23hP69v5w+/iWMGXEbIkWwzcFqx1Mo/IXA8U3s8vrvRT0gAFvrpgs7K9tPlZ/IhVXjMrMNGYotB5
jXrDKzeNN0uUyWJdtXq2e9dwiJ6rg5Prjt61O2GlXGABlFjGIR+twpgByj63LVPiUT2aj70+VxIb
yjNdzl9vd8OZWsKRnROxHknBihL0RB5s4ynj/AKXAZPRpdX1a4u7GA4kLTIWmLJyyOH0SDfNjdq2
3TWK8mhkfRAINAxy555WjTxD1yYu/N5X4kPgTCT1erpmTWPTtla7cjYY1j8OcNIZSd5Trgo4fabi
qvMyeFw9Nd5A1DHmJi7dS6WmZcTZxH8804BYMdw0jhQ6tuMHiEL6muL10CopGRt2uhCi8cabS1Nf
ywnmHQZAFbjAkfYT9IgcTlVKr5lskb3Z/1mHUq+OnAcN7DsvwiGOA8KsI1/lLvFs5vM3uWXnXHfe
b9icJqGthwIuj2fE45RMyxatoQO+wkloY9Yq9PHeAcg0nDh0qJLGGWrM9jY9Ld7+DT+M5dkmIlYN
w51u6Kptgbol/a9vY4s0rlP5aRfl3szBZmj3wnfzoDxqc+wCBWPmJb4niFr8kpS2xX6yogNJuRag
gFinRo/qyFbXWooLEPmIgtWd+uFxJ2k+Y6kqoI3CmMJzmtdGWxQHUvjen7Pqhg+Zwia2kiqjEb/M
Z3DPuCDQJcu97jpxs4u7fOP+kEKl5TZzywiNV15tfQW9vqrFhFczPLq6HZOnzgZLe7tUfgIFXtU8
8EWsjvL63aRPd2xsdOBnMXdNWJs6Gp+nVybWRzi0TpazmvMWDtg++agO0sG3J9goxz2ZzI3x/emw
PXc5nhOdIDXCNhehc2PhovMEjZheAccL9ZJHOAG6lysMIgwhjh8dgU4uvjXPD+t4xuwb77aLG/yq
LQr7sQCftVgZTD5nDIN6DO9gLCYzuVl3ejppbpz05GmT6fkqAaLtfP5ayoWzNyB0fvhgpws3ZA0E
0J93wvwwktMhAngQT1BGb+c0h73zPb8qTJQUVL9PhTFQ2esPS8zoqg9a2yVMuyluyKCkjlvom1LG
yaWYhVApv5GOtDYwhrHlxWs6IxGl7gmfgcUJdpJYqFmfhoWu2pr0PyKRnIErXGBVbdnD98XqSIwU
Auouytr/1D64C9fxPwb2XMkqZ5n32F/5+9PVD0PB/ue3oojPz5zj23CkLHJBqhdaHITK40FdV2jF
bRfONiKpdfk4wOxIm0+BdWYnPMGYpyq+46Q9vEniQWcZCI/GXYyr09kd0cNnHu1u0NEjjp921AeZ
Qqjgob/TGD5EJZBB0HRejUrHKUpmzZAOyfN5jB2if66V26ZMFoL8/fxg12nNdsT9yhiuNLR4U8yN
Crg7DbJ1XjCHvSPH1rzFJ69Q3IUuCGZz/hNeSiSPz+o8Fg/oR364Cpz/JhpKpIyFTt8ztFZPCRdc
t4WImzQfmuTciMoiFpuwY00B19Uxkclw7hG4IbSm1K0furGk39SCJZRe38nSgFHNZy8c+5xmlEsm
qfbNlOUOYxxS0y0T4HwhokpmBVH3DVRb10MxkucclMPXlxdefJD5X00PGpceacQxmPgIneP/d+Zb
3QE+fqrsrY/I7Z2/Ve0pVkQ+/TK6YMIZsCK6WU52r/je6IKi9Dy8iZAW4wEDuYUmVKvXTSWr8nr3
QHZvbArtuZXhiLPGFaudNqahVK5tMr47qRpu6V+wVlV0nGp+Fky2X0Rm/xWfCLtyU4z365iYMbLb
NJD1WjuADEUlT2MjhzXN3gcnZ/fkpCsOXBtWq4wxh5ODsQTBbqOmvDKRaLHk5jWfcMOJ+ldF1K/X
cbhVsDxi51X3f/EsLNhhRhVQy/rT4aJcQAUlettMzKHf84zu+09i6wOg60JRYnuQQteUTxvb4Sox
VIfvk31DzMr5ShX/zNy4Sfu1dbbgc6HuaEZPFKzkodFo4yfWCn68C0f/6Qhc2e3TvYrH4NOPxmgJ
Elm0+IzZHwtuDJZfFLameDlB5XGdLcKl7oW3To0DBMCVdIdTjp2O3FM879+08XOP7VCHMbBfiBL4
UJuFoTsNuX3vEYsmyr6l+I8dGJJF77JRhs3LFQCg2T2tlQnN+a2l6mYVitoRomYiexsxXcd4qomJ
za4TkIsk40Z7OKemrEQ4LpXsFL1FSko1Zt11v/ik0KciOO0T7hKnFPhDj1J1OHZJQt02NkOgTb8W
j7IBmY5x1QR7OL+Xua/OL+liPF/tKvCkvTMNjyAQgGAv1LvnVThLDgdgZemng9XopHa65HwfNYpy
9eOFuSuV7c0IwVZGG/y38BcfrN1uG9cr+kkmy6hwg5I8XNcylznHHoRWpHGj8ct2C4tfE9G1aOKg
au0mzxoGJFfrcbT2PfHdQxTc90v7Jt57ZXq52L4nK42icujPKOUfVVDYA5UYczvxO5ic7DQppoWF
dLlEZITQzhBPvBaWZ58aclvf1OTyC8+Toh+Z/QTaV9tL8KSU4p/Q+4Tzjz9/cZZEP6L02/lNoVee
N8EU1JL6ZQqJShwBzPTBrQcyApXa2m9ZxVWLaCpMo+23JUocDEb6C9Szx7MXFLZ0FOXvvMdnFPG4
rB2t22qB4RTiPWeHJQpNSo7egA5iRAIM/6QXTIwhG63NxWzBoEfQpa9YV28+n42NnnW+sSDcYKPF
voOKp2xjr/+jeGlCVB+6nRohv7WOlKr04VFdCgEjx+RLCyhniJTG4LBgwn9f99HmeyObw0H/QSaI
KJDevkFU2kx/DJzfGyM6G/G+Nxks2mVQWXXURtd0P35PdnsQWancrPC/KE5Vgkjr21glSTyksFoj
QqF0MRG/fjA1bo9zooESbLAWPQ5QHPtYxcMh/xfAX95AiVpNuNZV97vBZZ8ysxiMof0w07K/kopN
muq7S/i7gcn/KZ6J6MPlpZBmjrpVzTMRUXgjE7VFEP1eCymIvp+5WQuTFqO4ohyFz7jyaM9p5O0o
Ev+sXbNqk7ABfXx8zrY0bPSIW8sO8OJaGgNKDK4WQ5jhVT9gWZHa7xVnL8IQbd0RK9yN/uJkjPb8
daChDv8vwZJLpFPQvnvxIMvC6Xu0669Lr7B7epn4BuYSvuj3E8pyxm+lDQgE4wjDCll3C/Vt6lhz
khh8zrGsbZbn4M5hzO7qQ3K0wOr+uu1XBADYWJEZ+8mjTP3sls8bH8Itg9EiMsCJLoVN5lIsPuKj
/OncyooB4KXZFVcfhhjSvaTi4LLdKNCU6N0ngKEEWNJiECwfwd10a3h+CCatJeW+7KEDTryo5ufh
h8IMCpVnM8ytvUSodPhrT3+EpGbF9ct+xzAOtUYPQ8HUWtXKWcP/7HmUG7Y7Q1jfXtVFS+Vlip23
RP+EHpYuMtfLzyncU4NMzBhw2hQosGasv/WOiZcxrXONDQPAJkejSRHYe63NiyCgOLf0Miyh+IEd
yndWcj6Oc/R2V6/SX+RNQtSUqWvv3LMXevVYDz6f4qGv1twCrTxNliYBqZr9GmTxdXuRfFPhxoM+
Xk4ToadZ6UGUUvi8m0AKbHltdb9jFVGjK1KlNFFJAa3G8XjWf6MkWQW1gWPtoeixhu/IF1T+eo75
uqwH531wPviZj+ngfSt5hKMMwjVAOZK63nr9IurgDKzc2gURlRWiSUiFVDB3MVSIiK1eJJw8Mihw
unNIQi2Y5ZG9oSOUIHc84PiAOwWRuDJTw7GLsi4bAfwj8XZmVpNTMCyUfeG6qTGERlphQgt75hel
Qc4eqRbVkvTefvuD7M+ChsqiG4mrXi/2iUf7V97uwvrMacGkEKypszElEo6qGjJUlBjV1WKHShps
fGo6zPwWfMMf/s7ng7HOCRPKugZH9J28HnbRaVj1fneml8X6J0C06IHbumbGenhmB1H1Islecba6
2CYpe2pXpL03s8fuBs8sv/amiNL1sDTNT5LS0sv/wK8c45Sk1MFMBBPBVlNIZQnSy72YgNzPJewH
lGxGWxK0INZxmCqY21G3hSpbWJRdVNNq/mXmn1vfXhXtzn/TR3F17RNqUpBMf5NgCgBifyysyDoN
jLSyt+BZUhnGAT7cIn3ypxxF17KuEWG3/XO39t7+TQLuiSQDVnmQGOOqhk3S5uaPUNtBXEPHq1v6
G3lNcFOfxa81qo10SRmp+ufsGKxcqfWnh8p932tQLAuqYFu/VoTR+VD7Suyi7KLsPtmlJuN32wHv
ZYNkZxSnq8eEcRzalzFg5l+Psaxe1RibqwGt/azZwcDRew8gT4+vv6M8alRoSX3va+ClLooMXkWp
p8p7oegpRiD+wB0G5S69Nhw69m0itjco2dW1q/xp0At10QYBMH7jOlXaySRsL0i+opMXGULEJpM/
mJDdN6xbg4NGR8F8+Qx/akHptdUQoDSpJWS3VNt6hEiq8JYKtBNpFoKcUXMDFOYV2aEPzihNhT+w
QjkWzZifIsW9FaucS2v41UDJkeepQtCE67fQkveI/H5StDbwl54LHPahl7LHIjzq9Tx3TGVYFmrD
FYItgrT/X1bjyHjmZLwMocBIQlwUVB4ym9hj+8fpQqpG0sKgY2I6NNDprBJv5hTiTomo+zjNG8CY
jeSnN5d2snsguG6tdzZEvP9rUqfjasDq7/EuPAtwVfDKb7+PJXhKq+L5cBGqcVnqKVijys2X9skP
s14DLud/BtB/sXo9K8Vsd/5PNRfjzVdKpGAoymYPpIMSR5hDGa2RaC38Lz/ICuCbVBW3Bf2Ier/4
ib1sJuXmqo1Kst2Cwv9AO8iZ/honCCJxuo75hq9fScDs/GlGY/0jp2MF+SZvG4BxckuV9tRtFbex
Dnihr9OrY95/cBoCQFpdcX5enN58hJz2k8PiKlHDmwTOdyee8bfYId+qdDlQda1yf4gdNoQo3Vm3
aArfqJBrvarY+JGqpufYoPzjfjER5VKZ1+G0mDsL+VJXuKTlk3XHvV+kL1PeCCgLdLSw8SDsrwiS
TlDz1sklU/xjpr0Il73IrSSDvBqxyfjh3Y/k0Q0VRUa5gnAuipHoFFGThYMeHZnYOyFIgxNiqETJ
MqxlyX9j63fJ2DysRsGTBGYkABnAqsWIjuW9w3wK4Pfyyxsc2XI80yVD8J8a9wIDoUG17QAyL077
LViKzJxufzZsoxOiex8TjsCZpIU2yGg20U/hsaMpxihC6NCFszv39Sv4WGTBbfbe5wRqLjVSJP3L
kpaGhiJ06NW8MciCNHZXQugBAeLRjq598Pds9t1CeQJuK9ahoKCGuaBQ/9ScXuSfuIjHy1zLEZY5
oq2E+pe3MAu7GpGaoXWXZv1/FFRl0HA5FO0G67NaE76kogIsDpbPwWO3rVIh8x4BGDZvWh6JvaRd
di6EXft9scRpici7CYSr+1CEMBqRvhEmo4y1Ay3IVK7Bbe1A/KxOCH5DxevOuCbCwnihGDYoBwrq
8IvJmxnjcLqIiHWtVGOd3XZmLxo2KGdXOyyEa8JKJ33OLwmMlWwWJEF1pBhZ14/UhCOcBa5p6El/
e8al+ZW5Ea0ivzKX4e0X5NY6KZwOHpsDBzRQTp7YBSKtKzTaSHXbsurHWOlrBMTK+w8YZ4QctAUK
SEo9Vlt04mnxrwCtUzGwcIP8vjhwr/FExy8JrAqsdBf6p0EIc3PhWc3yRuVq3U/kJXKT4CGhhEvJ
bfGArthIIQPXDMXjp6ehgoE3LggumEa5rHw3fiL/LUJjCBz7ECXxavnwTUf9Lgkph/ifwZG4nfod
7WyXQL+FdfogDQzmeHjFbwrULk9FyItw6pEqVSax7F0nzdIu6R8h8Y1htIcRv5jFHWxG/jSUnDJQ
JEZkhDN8vgkDxO8nBTgJSpLGcpSg7aN2uw5tr5hZuCBM7PSnlR/FJR7tZfxua+mNKDRWbBtYyIhU
2Q5lpSta/VU7PYAQfZd55bi+Jnzq3tmBz28xO2GyEI/eBjd+Y5/Cv6sVVJ15ZwKfXJDNLv8WbNOq
T4JDYg0JhZy7T/Q5+Vy5Cfqye2Eq8YG4rz56JyUtXLZp3oGq57nKqGIUV6LorJ8WtKYCNkD3Coak
hjxktV+IBdFRO9lACBBKYoe1G/w8kaKRK2qRhWXq6QxIu8hIUyzRjt+Zjq4dlvs5bhZMtI05UYU/
25MxI6vleHjkemXUbMPml5Fpadlb6/Wrm4MOhSnPOt4lNQX9xpxmICSp60EejCWWnQJkDJDeGyJ1
/p/NKsYVS7lFiusv2zYAVMfjZZAV3AQQ85QfJ6bDRgkVu6X4abBciR5NZ4DDed5srlS+gLCfhU/p
Z2sPMO1ZwO8WbhV39N4PeEAblf+VI3nyJQDSadAPmTXWyb19hWLBj+olrhcd4WreyjqeMkQUi32f
vEXUZtHoSsGIgKIymSMgZVQQQzhKX5aYgiGChwb18110UAbNqEOIsbooV/NDW4bCaBxFr84vwLUi
ajbDZ9EFLJ5yO2wVtGKqIf1MM8OLTnRzKihaGCEYJNEAocKEM8u3DOVXc6yAUeLXI358Vtre2ObW
HcbPeqXqUwpQfZ5pMMm76rQONnztO4caVLxC0wApo22x8Jj1h4Pv/Ci44QjnBmhiA46jNwP8w4eI
yuSL+MmfyJ93kYglF/ARUwoq8Wz9HIyqJ5L44AV+pkq7osW6XSDxOGjPmy0FqCIORajHvJTE44m1
p0PCcntSRpkPY6WlkLw63Ae8NWN2npJusIvEJ67xS7i2qR+ffyNMHHeI++1x19EtV9hsMT+Ej0E4
0OO2hRaOaTjDYZ/X6I3atBu8iG3DuG3/hUNvgr4w3f+Ff1HPoi26S16bjB+BxRP6K9NK7Y26O+Sp
O0lyuAjK9YH67tSTLFf8La2gOJkBXoQdnIlOx6uiefZwi2hcWerneReIkC6mgbTAAcQZRoLzIG1I
ZrhZ/I3j5UQV9ivsLqOw5cTuugz9KjYY0p5gYWwWXRSTd3NhgdAUd4b+QB+KRJ4VX/RAcqeUr08I
Ghia4AsFGj80VSSmULkQ9U9uRJDXwYtSyZW9bOLX7BL39MFKbnQ7aYMKRHFvbIEdAhqNisWogOSx
vQJBNJYxV8cdue3kLoL6WdFLUht/BRiulDEDSMhNutggcpd+q6lHzjxkOD5i8HabIh0mzqXR9gtv
085rOpoZkVHeMF7EYIkCHnI5FqUZEvBWdGTk4Afnvywi3n14VizRhJPLrFutuY7KfGJMW2HuXOYe
ylvuyaIP3YZQDkVOka2xqHhaSncmfa6BPBJG6rBDi6ko3V9iJ3hqV1yNXmsEOFeuMRnxVyD180TI
/M+tXNH/npEkSJ2zsSfC4SUJIcASNmQxJnm5r/j0pYTsWKwQ5Ie7gpP3G6g5HcENcAaQ++G3drbW
9FjwXXp1IjoAkjzPJul+xJt5qzLa0ugTzPbSSitBpSMK3siMjZXW9FY1AuToMgVvB1bs7IgecQ+8
jQ8GgmUFp5cpwlr4/e3Sh5GvrYNebDF0ZGRRFNqhbPCnH5bDkcbwhXomuPnUSAFF6EJstacU3YOE
qoEOoseuKfqUtBL8egaf4piYbZUaspvcHiMBbs4PRoHAbrb2sfYXVvyzF9tBi9BcfXZZ+Gsy53z9
RewgL8jmj/dtcslKCXaOOmA/nshkbHRM3jio8JX+OUjgJn2hloEAuoUxfglr4mu68mms+JS/EA1S
t5AGyUOHlygFSfXlMVklDHm5Kozl+PCTK0epM62fb2LXbV9XhgAw6FNtsmW4P/ELHysLs4W2oqc6
PGMPojyf6fI1kLI71IcCO9ey0jr8L/mDOop4mwVl7sAB0fYBFMTGGzNx7UlsSQpLz9lCVA61YVYJ
jSJbNvUVo75g/Cj8Kozipy6FGLCdTuRM6wsFGBCCcvkap6XQV6+2dUtS3+53yyGyjhpVYsq8ZdX4
hTHops2xGhmVMg/pVnvwFgkjFIIiu5gnIyDRGLHqE7d1FIYISk6XkUW+nEszTJaDT0Em0s9DqJTw
FFFKEbdjnhjbbNRRMxafyIvPnT/t58qHPYUqJ4I/dV46K5UukCMP14m6QiIOu55yJe8AisaiJ+Qs
MpdTker3Jr66j0SZGMRVib/jfMwgl0UEgSxI2Zn7nXvlIrWCsCoog/D7AISLH8Luphez49fkpen4
ytAfbXm7mDStqadBXiVPQ/+WQ4qEUmC44oYo5XSHucuZeEHX+Q1NtYYVUdXyAbINhdHttTyaUp3A
pXVZWrk8tWdTlSgUPMgHpM/io/f3lY4NXaNXrOEBXO/hzMLyxt6bYFLZ9RqgpreKPVCCz8+MipN0
pBSd8KKTxR9HK7eTWIilVsfYrjU3h4I0maTYjL4Xk6PoSeEewpglk0z8KhipiPusVhueN4I6pTMG
EKsyY6Bd9CC3cwhCVULldTRB4KpGq3vYqEbf6P6YcWInqOSWPWnfol7Sl+Uvo2XUdUvczHeu9IVZ
COdrMiGgrOZBdyemWNwInurgv0dR4rjbzC3ja96t+4ShGDKSSeuxWhebEIIXAlK7twpclruWNGZs
Qb2xlgT2Y9rkfQ2dpmZYJ4SA3UcaAafGAtfuOWOJLi3xwx8MsV2/QvI5+JYOT+M9um+XNm5Ze715
xBATDufLZ9aNPpPWeYIsKwa7wl3NRSY6Xdpb86OOd+0+T+mgffU2GF9QeXnIzubvzXefRfwGJ7Z4
J+8FHCAsR6rxeYa9hO13GgEbIMhMxJxP5mM0YhxhespC/oYF0UXRHnfJ/AGcK6CrPSAR6cSZMVe5
LkdKmLscv9cyzAe6RPDQ15fCLaj3iYo2L9+MsW9mmy5GOp+tXzv88wiTPWy15quTE8ElymmuUDIy
2McXoEiuVuTsf8hPSuh9gB6ZRER4x3FRk3MSyajVPaHIPVJdz0ochS1mQRp1cnQq4S43g9W/091V
ZWNpd9tXif4qLpYMuLvnXQKOBWJwteSxupmDpL+GFPFsBdEBHqQj7NLsB46oR1quHw4D1STvuU2R
woxEO3l+s5omBThTRSMuAuRQjKF6HlR9Hn/r7588wyDSrN7/PhU8kMHj5jvZfYukyZC0Xp8ENjPn
412q+yGLRl8XAu9SAJuSQ9ZxAR+/jVSBUpwU0VDE4zkJkkLjMuX4P+ocu1ZAOfCqB2ThvRi1ZRc9
NK7mBhSgecpMsgIm1jNAdtNUneYjbiStR0vnuQCyVgXl4jnfQIkVmvGpdm9xzUUirzsjvVnu2dfC
gs/8gGl/uTYkA6Qi3lmuZe3oE1zbg/ng3jz7GuoXb7Hsno74qZny0XY8m1+fDYqeyjYZiXPLkf12
OvgN/QraGDCcPhuU2nI0WMmaksR+72WrHIAYxZoxLXZlzi1rUOozOctbsoiY4xB73iPEbDuzP1C/
kRY8CEMqYXPz/YIbvlUHQqQxrNlowsp5XKkddvb6+lzClqxVvEJUaxVPxYlbiytuZDw6V1TeWl9U
1Hjj/lEU+VF/nSMINx74w5GtcGwCuZzTsib/RUt2CLxCZAYT2ks14OFVXIJPuQ4EMP6PaLSCsKHS
CWfkQyE/ZY/Sx/xwq3VqtABApFWQueIMNEGcFNDliknC9Mt4OeUieyvh6HqRl+ehEgO+jeKm7vd6
VPqj2fO6lo8yg4OsOmadSNIoK3xa53hP5Pfn4W1TZE+COxaDTZfbRudXb0Jy5awG4CBb9t0dOAsy
upKK1HNxY46uFlGlcaZw6zFaJUqRFDIAZ4468iTUiu5B4liTs2uPZy4Yyktf8vgQjHneCj7m+zcl
/6jTisw9OPczzkh9Zqi8n2fyyH1gTFGCl+cLRz67+nzNhgybgSHNCA+w7ZF6xZLhDvkRKl4JKp3U
J9yvJf6lx+y5oxPbx5E6zOZwZcFX52YhoXsvvWHcvjsEQH4k4zHnlqRQ1EovDL2O55YnI7nuEqAT
ZloW7y7jny0GQo2GDCBfmFlvjV82tvwwP+eKzdK3cIyNF+1IGj5446ktFqkEbuZrH4l6agxn1QSS
bc0A+0QElyDEU1CbHF/C/1hX6DA7ojC9Qm4kGwAU9UlJSrTtbIAPjKTILKCJgYTg9wgLtwCFQ8yQ
Ifabxkbvlbzd63KLnxhfeAJbvtbiWZ8amiZ9l44qpAS7xUpnZq40P/I2tdnt1dayj5MwFGsXbWB1
N91U9XuMX5b97uhbHq9ErI0rL4VIeVrgqRK+paRXxo5kFoUOf1sYha3/7iwo65owkfQvDBChgczw
aaGfZEd2JyCY6Roxt9GLuIrCxWSWsKD9loMz9G/7wfJUumeYgB9tQKwTOURBZWKd2A9KrY0i19RQ
2uQWdC7Ra+PKtKDq/4HGbvNAJXaU8zD36A6c4mBHgMyQqEwj9+tsH8sVWrboJRkYiIhU7FuR+T3b
TT/klgHoEDDfHtwcuiVMjIhFjbllWZBgZD/ZoCiC683sH6eOqiclM5Xdfk8EcJs+a5cjlNv2xIsy
brS6C5kcd8WYFNDNLRTbkVIRFApCb17NgRiVhKcOmTASqG2+5DQuyvVopqznaDCipiixVy6c0eOu
E0bygcsQwqGgjaUaemh2QIJcd/X7TaluZfT3CJSynOYo+OsUJprfTGV0eDMeDJr7AJI9JQlm4AFt
AnFnjyzE/iKUO8tSFIFNLxrBR6bOUldFhcHO2LksdaW0kuntgecTVdw/zieNKhI/qKFoiZuuNgIU
VLUBOjXf5jEnPDec7Rpk4I3QFaaZMDSL0t8M2RcDTs7zMJRNgIfVkgg1jeVV6LP67goBxzrhn87N
ucRu0jglejuSlKEkJc5CfFo8hCc+xKmnuf7sbuE7lVJHLAAs4+mYhcTpR8rjJkZxAWSaBSoo0nEk
OmiD/Afl6sdfFJKMCsgTM1Xg9C4yehC9N/xUNfTaPFviRycHnhvqN3un1JePfNfH7xlJHRA553Mj
xFtXaO3yxrZEQ8o+4piwhfJl/dGN9t6BVp1v6tFZXzoxGs2UsSi/RX7za97FSK1D+bKzLe3EEWkl
6jErhNPJqsfFKkpk+9OaK5TK2dGMn4eIwiaJEZc5ywZpT/zjOfotgQayf0tcf93wqyrLpQ1Xg1Un
Fpqd+k3gnrwKhmPsEkTDmcKw0TP7qYG+9VCdN5mRHAcS0aELz+34UOdwngjjwrQAmB36+4vn4+19
mxe+9QzKEhBqDoxNvY1WtNzityl5c88QfRL3MiGSPS39Y0mm0Fk5fAE9EQ0SzQb0VkhWH2C0PFp1
FtRKyDZC+ZutaeE+ZpUuLeV9cXbOd46mDGiZVwhY8OzqoL+/c6w+QcPm9kpWo4HE5j29d+KcAtmE
xyms+1hBZKlM4cUpQtpsGO/JUk/xvMc/RT+RlEX3Ykrr+CLIy7NNyYQxow7s5NfQ4yFF/T8nCkZ7
t/y+fbaouMDKDmtHK/FsTiF9JkEJC62K2XI/jhXT7BfUTPMgT3HYnOATmkpkgKsuqtgyqn7b8k7n
8Cj7axJR5xfozTz2/kQN4VuuBuVMB9b4bpPgIfHzpKEYDRps1c/ofXlwwbbtqmFqgzO4E/RYUCdu
qOvJYAkD+eOjQ75QuKeYRRxCQ2MZLswGg16g2jyozjybVcXS979pVM2zUiiBzmh48W5VIyVpMztK
jgUtm0ceSA+LOsku/GAGi+W091vA4QE83C9m0Mz8y5g9QRFG97B4PcvgA5Uma4IXXpJOgO/fbro0
5TkhrNsiN/ZEOy36Nn2LkjhVUkKRDHUYSC+4b1b51Pd/eVugg0rqKLqVB8Bx9ujS6v0H98POsGq/
Lygqeo0l5vVgIVu4fw8Zs4gKhEjmXQl5Od3dJpKxPiKqQAghKLnoc7TE2/yfRMy0MD3+TnqV4edu
KnARjCSThjzk2qaxa7ACXp9rCvzw1U0BldL4RO06cbzAP5LyF4h0KwSWAOtQm5cdjiHgSfGUolKK
eOfVzEXDW/F7NMIkRaLBI1dijMYrojTFUv/HmqQwg9L6t8CDIwJa58f4a/HF8y5Xeam4X+B5gzH6
cXPWlehndSqP8KP68kU0RaUEt8vwjtMUhYUs7cofBBbX1imMtOJlR81O20ZEETL0WWxflFOp4DGz
MMkPDcUNqs5+F8vvMbsO/NHTTPgP04DEFrUQdXwFuRwE3tAWuzAq6RWfcJ4+XEOwAt9Q1/QTOrKB
ZmDJtcOk2sudjcJcpI271S4A9j6/mDVyCPFV750XQIRnVaYVMm/FztLtMtmJvStt6pp1kA0qaeBh
Ox+d47uWTAc18RBB0SqRL+m1gjcp1S+abJTmWC3DWw2uanPdSqNU38hBu/kljRIBvMgpfRkPOaIF
DHE2IVBV4QSjL/wu2A08gVce17ki++x6MtCpts20ITTF6OnO5B22SFG3zdKqUySHhH4810JdkX4x
fClTCQdsl87rvcfxr53H0HAsnbSX5uNH+is+jLrgtkTwFCShmxY7GL76KRKEua0TAtGYdVzxwPCK
K9NEBhe/OvRM1xfCl3vpAqk212+kTNI4qaXeLHsU38RXCL2OrHCthkC+zd79k7hcHuXKSmEIkHWD
IOml1yhnP3R5/KreybnkMb2vQi/FgRh/iiHz+HvteMoZ/fl+y83K0yne5MmmXQ6uHbg0muGYwUvM
pLxPhIdz6WXyAHmIqJxjU1OwwX/KnUpFE3x2Cn1q+QxZ79gjlEqmmNcQwupgD+cGjowUOENHpgXs
wcI8CIR3yV8hL4KWbj3bSZX95mz7iAGEeoAbpNWAzD1SGtpmG/9J36yRitlvTQiX04ySknWeZJrO
lM1stglpLJ9l41r6tExCd2DLGQpQEJrflq2QUvtyrmxYpjvV+GiWqYGA0i2uhAxQvJ3vkFarZG4r
4FwsHIFlbKuxXa7BL4UMzVccoAVHrozm3s/gLh3LE4zU0oGIt3bs4Fs+tn1gixZ11A4+nOoFHbnh
SvsxW569iCjc25nvh55qmviCqqxMs1by/EQeUMcwwXTUoCzaEzuvgqIHQiPXBboHEuA7JdEV0y7u
Aw0siUA/K/MkHA+fxsCVJ02vx7iM4FhjyUvaM0xnN18bSinnNqoI1HmPPF9YmwajZ+W0NxR3/V3H
kWTc40AAf/TqbQODnqQsKTvdIO29nWvCJXc2kpiwOaPZmldvPWmoXNKOGsExu5KNhsG6kvg/ZEM/
eiHeHyAOiz9NvQyfk1lSy7VBj/zrlF7DN4cF2XXsNww0JdMdWnP/EPyAnJDxLtaa1zW/YS0cGLZe
ebTY20UYjVRTpLYDEB2I5SdTpiwLSGT55qOt9Yz7HTzBxhd5/H0+grOA0m5skV5SKjKHbOYpinX9
G2OKR8i9EwPgSP6Ew5hBaCN8sVLvFiXdfxNi2r/RFObNIXyftVkNbR+tCkPovhbn/c7+KqWdFbMV
zMt2bCQtNArjoCRJtzqa53SisE1nLf9BHwLgL9M6/qF4ndaLtKj8DfZ54MBgG96A4l867S8eXwac
rq6bw7n7HGZksy7iN86w2D4UCDbFAUfmfv+myAHWf5SY7iDQIIYKvnRQ9/wqcWBGE9cHUtKWJrRI
lbRkUh0Y4/WOOJeufw24lgDlcJZTv7tLROiNb6w1F4I8XInLufB9mfoWsCyrZ0vOM2v0etFz0k3C
qzNc7Z8jEpvjInIAUdYQ5TSdDK6RthDKPJbX+vYRb9z+b7/UaEMZD84DSBUkAHKPSrU3K2we5yJB
VlHWVDaa6EXz4n+bu9vlXCZAj5MOeq0cCP9PfW1wwLuNR1vW1yY6Y2b3yctsTeK1mBLblaMklbal
Rqj407weKoB1UIzm6fkWOdrAJrlZgqzHASiPIUAzc3j5hUliFah7XyjlrIIqmWlyuYOwjrrSUS1M
YbrUwNU2n6DQwQEDVcKffRu6sd3B87ItWXBxq7ukqzge4w8u4+lCqPHXPuW/Ll1/xH7zoOKYAan8
6kAprN67I9R99eO6EaTRNEHy+AgWcIoJTOLE2IPERV01KcOLQCYi4wROlS19gfC0fE7L7laBFtFr
a33R1Ut6ktp2yALjfAeOGD1XMdhMZisnxiy2HA/vhd5uuC2UEHXEy7BojYvwqV7Elaji8Qtf1bxr
csYqXMJRHkGm/58dbgf16ttqlu/xnsIdrBxXImRhcx7YYWoHS97HHaIKhHFp2XYVGFwqOTdqpHo+
qqAGfPe9U91UoZn0519s9FEzdX8T9uKNlbSxMUxZ6wmNWeB+xcd454z72E/2V6GngzB/9AoZZSkj
UShMsIBm56rKXQvjX/UXqEMAEewNeDyr0KcMAO7X4P/2HeD1+YZ3x/SBTye+3lXTy3kAzYkC4+N6
efWJK3rsOte9lP11Gqf4RDYhLa4DhBiwQIYixv+FzDx0+IZ2hLbGv/uc3ueW1ah1uG0Pj/wI2LT8
073/YOfa1aLPt2BR4yEjX0PAmX01LimfZ9Vvbe7of275pl5LQ5tpJW7BFZ3YBoJ3tPetDbOWWWQc
Ur4FlpdvsYMNiQ0h7Fo+GT/NHUnyA1xwB4ucDBfpriA9+yAsb9opDpH4S5ADDEkI0iR7HNyalYwc
jxaVNtLpcmt9cuX0YepAvUJzToq0UmQBHzqbVff1oA2NJ0knFDVrGvlkKOP6h5FltUs3HTr6Xxj2
/KY7KRIxNmhOHHoLIQHYc0orrnPTQZWF9la570Cij15EN7SbYkc8BhORvvMs6uWjbo826ozhyQV4
ZW84dbobw/2kekFepi1hy4jX27CHBtaukuUFOAhc1q7jjo3nQudQrQ+XQU8wLfg7gNcI+1fZ3/DB
On7pxDyk6h7rvE0j9pPUz60VZcaBxOhAtknP0PJVHrcePqPz5JmGmpKrqb+CTnTahYqjalJ8ZisJ
iztk99ssxEav8EWU8U9luBoLXyngBzL9Ms0YijAirfu7g6M9rEbiHNfBkOoS6VP3/mPevBW0EWx7
cb8ozY/Yustk5cD9CMeSRkIFv44chUx64uAAUDjUZs0F6B4bV3zp7pXWbvx4bv5zR7mYRX2fEUZZ
opSN0E9hQFgphYy/oFmts/JDLVnmATItzmGMhi5erX17HclYvlricuv+XtvnmBwV/XED7O8wFX5+
nH44zD0jatjcSRk3st+q8GZktncEwcsqTmtAhpNdxonAyOpjVMHiT+55U2cvMkGJhfZYIK5UHF1m
fgOSPoXt24nSk2erFi0gMUUD7JPT8T6iZbZY6oSHq7369ZiVsShdM2Hiur9eM9g23t5RnTR3nnmJ
N42tR+4I7consyoF0rIvleNzPI7Qy0uomUZqsX+26hY/eNIFPXKxCudqNoOLVXxxcweEsLNR/6LX
uC4z+jwJsasxKfVTbL8pUcDPeC3ZJFhAdLVK7f0nx6o3DxzWnIraB0fa56l9rdnN3bp3GYTKthSX
Vt44ElwgvE4yNPfxFD+Tm0lk/+Sjwsns3Pz3A8Nv2PZ4YXaJsZWEU/kTcJ55ViYYzKFaF33hMA2w
+WcwEZvUCRnEUCA1f5YFFIz4EjrctDtgzN8hxpzvdaYXn+LH0M2VMGDDPAoadHhYSQnKMOfJU5V+
VegpJEb2oe/iL6svraeUskXeDKBxQhm2IGeXJ7cpYCCisNW3+FbfTLuyyL9blYAbVyWDMGFbmShK
ajJCmTXz8o3bRXgGs2TGM4Fr/yi0DSYhlPAdOhWUnDD+pKpXo5RnGfshBbQnv1cac7tuqNFHZol5
cXmyik3bWz8+fAYuh71kavWqGd71vLQjBAdKR8sLrPhOBHFQEHxKkJiTZrTjqPr8fwy7DopbXVc6
xZfWr+otvzE9diVanmWq+4KK86bcC3EizXIMbigo4EUBT9KW7SYU7u4wDfqeSf78htVGtbzwHmSD
bHe/M8mw/0UvLs1UiPxolF0ZdKFEofmGm+pobCK2NOyEh1A4LC5DJP+c9yKSg4wTO9KZDYQ7riaI
qUUhtEMh7SOIhKyO3ZSfq8kII4wLIfG4vwmHnjnPcUe3cwETsELHd6hGdZv8EFEgtvENu9gxqYBa
bD9sxxz1VcS5joqLGTcvRSumSqvDFKmAg7n76IQ4H9pnZ/Gtf5yPzi66bvYAK0XDoLV6hZnqJsnP
xJUy8JtJLa1IxO3Q/45faWh72NyHZygfxhoRljSEP2tK7Rb3Wjq9zLg+WUT0HLcS3J8R2QYaagaH
NwBQn0xIN2eH6nCfOPREZ/6kpK+3JDvftobeBqU97zDVD0AqUuuHvaj4JKfk0eQ+sOkQO3u+YmDC
ZKV9S2kHAThPTNYkNAXgM1+uYISS6s6upHkv6rlweMsrFP0AaIrpcgFUwA9rMdjxSn0Yrli/sr1b
R0IgGGbowaJ6ShG1HYZF7j8VMuiyQ0mNaWh0AorLucnKIho/caHNuDPTXApXH05i3iwfVe/XyGZb
gVxBi1UnVb8HFs6T0fJ0774fKMU8F0KQDcD5/+qp0Ricec0TtAFmZyVrPKIsg++QFeIRrxJk3L7L
+8ezuXV1rn3lkZuX6DH/fTvUvd8CqLpQFvatensrXXx3wYnhCYPrkJ8CNjl0xIrlk/cYpGVooHD1
G4kBYExBL+en/NR0BE57R1RVM09OPGRSRKY8asBficbJMLGAtl/z0JHXlwMHqE1XsMed0g0UeDsZ
jGEwXGSRGvBYGWDKd5oQuch2x/qVf91kA9XCBQ85u3MN8PGNz4yNqeJTEa07y2LLN1AOUJUAlAbP
Mpp5oEUHmS4BXcsHO+CPSqkoS4av/nLwX605Ngd84x9RzTjnaYtBOI8Qs2rspmXqBU0DWcjnWWUF
Vk8ZRLh0todIl/94lEPX38ubD4uqYT/5WPZGmaxMqmSdbsuY9dDzx0xsvXhuyBHlGFcJXvhk7r7v
auDFk2yTqXfb6Tl8Rm4iJWaOD68RQ09Hw8ByApEQdr6ohIz90X5xRcRpOO5686ZH63y39VyqUodb
faeSnD9lVO8olOcoatcSDupJk8eXZyg11yNLqXfRg5EvdQbjQPMj9GtrHp+bLfdOTIzitbBD+sqB
9LTbnGiTB9T2CJgkWLyAiRtF315ZwrVSRFjv4XG3EXg0RtmNUfoGthzKtsSmUNudgVuWu+X5bNC+
mhJZATth/r3I+EwG01IsXd+QfMERSARmX2i05tGQnzg4qQ1d6Fg17fiPUsXteTeR6FTWHnx1hk8s
r9VIJn0/wf6C3KOtIN9Zwasv4NbDZwvali1hbsiuMuK3FdHJB7mFOCUoE5trOTbeLid323f5IdBR
dEkKLWCYodi4hn32WDPeMETu92Lh5QFFJHpQ6r5xzTggjCX+5xQFNR/L6W6Ex4SkIX4ew+meKErD
etnfqfmpifaL3pWXYBCnmootVwTAm80ayiWjQRflsc98A/5YUwTyBF0zjP6ou4aAtlNNzfN43zD7
NyRdKkSMZe5luJhAt9OdKVI3Fg0wzkI/dGZZv0XvF4k7HTKlqTsxJdzRDjPPH2bfyEzGqsGqNNvt
q1kiqWqEmdDKxBEGLdEz1TeicRO/kSO+tvON+Z8HZ9ki3ibQoNRn5gC8StrXWK+EQmY06YqgJG2N
ueMF5WkQY3GOwIQhME3MP63mtQVztv4JuNl4O+dojAuvagMDqPStMRF9Xdr5698gvo9Tmcmvujzj
a7vJGrV3rO1EWHYDe8cUwSe1wm9iMRUXwqp43nEZm/hX+btITb3IwcR7HkXmZD16nfy2DO28UnE4
3sYFmKpaJvBMhxnp57OMXnxGmT2mqY3sYYITRqvT7Alc6EjuTyPiQhYh/SPuKdGJrOVKxnVa0wNg
G0RdOioMK4KTzrWwzHXIRAuDpzK7IIC6HG0e/7g4utdAQqscS2HQ7hOFEExHBCfn7OTPSllG5+La
sB5Zd2B9dAwH2iNFUlzAg1TGpavoFyInf5+yER98iZMCB16wW95JARPRcDpZaRugCelSIuIbGdYE
IrjVogkmmGh8KVz0inszMYDwSmMX5MwJLofjrbLHcC6PXiQ7hW3J3Qo1xK+v8Kmp+qFgtPu37oZh
nr9GQFJFTIQ1OUtEgVIKTAtMtStsPAYbxqtf79DgCF6rGf/CwFBzDUeJiR56ZucieRc3v1Hn8+oG
vJFX8JgQ1db92UM174VMGY4MVa5KvUOU/oZ47zesDovxcnZfr5UVKGK9hjfe4LFbezECYyTbUqEj
HeMpdbTHEj+Td0R0kye0p3tECL5VAFJF6kwC4g7y5vS8bJayybalktinkFFhvuBdNymJZTec1O23
2rPTaS/KrL6VObKzTtedBq37E9sL+Bp/j3IBHX0S1iieBdhpdZezGQm5AUjeKxkmNzGAh83Zd0b7
2gGY20C71YZ/rQruXT+GnZpW0nmemyBqPJEDdGvSvbeARm/7Gjt++Gh5++hztCxrW4ADDZjDB5Id
DihQrB5mr5xnueVxaK8g8PbdCiqaI7xf78d1i0GU1Ujj/1cHytbWnT93CfHES3NnyZZe3/PTXEkX
KfhXX19xYWZS4qmSLIZcEKRNAEF4gMVUHZVU8aRIBd5/SIyCDlt7S47UpIF7Egi8Z/DDM7YZKFHE
Id23/z7cq/yOzzUdt/tjjhzSN5nUrNsL9VelRfaD3RR4+e8GvADpsDCbU9eWTlbASzDuGT/juJ2Z
SbveJcSFy4F5DDcoMGfSSUnTIOV1iYKJWIX5CazRpswUQVM2qj+OSHtseYLiIrfYiUXmWhNJMGxl
QI8B/V2jW7oAqci7ojSrIxayQxI0Tnt/ihFLhOE5B6NISxFlrjwNzotNVM0u805wPcCwC5iLk3ri
lttqFar/TLsDbHV4vMyXVUO9R8WYQTDRcV4Y5l1NUZ6DKxc0PCSfAoY0GWvAW14FHSOm1tDmhBTx
yKrfq8Xs23NcTYIDgsLpOwLbqwex6FtO0E8wpvvoXdyvltWvl2uGNrhafoBQBdFQPvkk3++LFDAa
IeyAm4AGnG09dCVjZ9fsgK2tjlpMoupi0SqyF2al4wNm8pxULV2mxmKeIHfIuVsQH2CWI3NUaftD
YVnT8gc46RF5hCCtD7dOkh9To9aNrM0TNsu6IJeXjb2KObXp/hmdKHy+lkr0F+c8uBzEdtS8J/p5
3Lltsc/lpkeVVO2WLN7aY5Li8WXRQIE6Ff6isjjG26C50TwEFCSfnzWwnvsjbVHzLk+1/29BhbBn
Mr1pwfLkLIhXrEJjGxiRzUVj0BksaXFx+ZSyiVqZncwpg1UXnrZxqzjrbBpOJN+DeeoxAwBoC2Bv
8YL15doI7lx14yUZSgDsxUT36fQMfWq8OveQMZMN92MLEgCmHtFbDv8azZ4l2QTBS6OhOzbPz+p0
UlcH6Lm2ozQ6LdXnqQKzMj29KC98FxwB6jn3bc2kc4OFIiEvhgLuviR/e/W33jkcC/vMFUwFAzir
WJHyizPpgWtok/IhAbM4c6vqT3nIPcX2mRBOYuo92gnqHfslRrbpNdLYKjV19KVNKBW2PY42+Ak9
yvmumMS132Y59XXDXBxoW07u9uMpQtYvRFS0VL662orDdNiMcnZHn9oaexmiGInh4fsmUM6hwd25
vJ+4wVS+lK34azqIenGlOcGqSpu0OE/JrL8vnqZALT0+Tv4PPNBp8s5mhNY625O2lA1WGaLUECgo
wTeocqY4QLPzbjUpwVMsePEk/7xxl9DnZSeIuez9XQtkhmEalwomESvFh5ybzt/F0yBVtqEfRtV1
ekyAeQDLpzZnEiuURNYrJjqtuUbNR2WV1TUvNCxkaLzcgPGOWSr/fDiI9NsfhnpF9sr9O3ldGBht
2M9U3DEu4Hg7526yHP0WhZ8UtQIqEK2bGE8FpvYEThKwjPgwWVbkZOFe5kzF80Bj146kw/pQ97fO
ONeLAUBLnVCg/CekiaodmqMMJeLF3RBuWEK2SZjBtyAxOM8RLbkve1H8SHinseXLOz4JKxryoO0P
6F9Bwyf7XXjaKgJadyQGg7dv8DkUNBbfzvGkSsBndAxO8pEyplZSNdt7/mHJa1SzxRRhqfn1WFtN
mZcyxUc1Vu5AXcUXuv9zDN9W4EFrn4yPxAsUbH+Qp5x21YIAXJfuTf+vrjfNEJl/cloMkA3h+JN9
j0KgXHmdtBTDjqQKqi/aOf7Fz90yx14OBCDp23AWzWX08n5Vl7RWfXpNI7rfXhspoglQ9V/1bVi+
c8THW5PqCZSCeal81qW8jgx/WkeE/m41r0XtdGpn7dIJlZwQMZ0gFGyHehSudAoCalXdc8cavek1
WKwDqWjJxwXshP05nuVtwCCcGCHTxkzJGBMFaDwqhAYCCdRoSfN/H8SSC9lRrAQWmXKPwUnQawOp
t5yEG4DaIYMen5gDt8JPBW1capnz+qcuQpYdqGyZ8OGd7iZ6e4FrvEesk8a9sqAPWKY/q0MmPIZ8
5bQbYC34hq2JWtJ8RPDl4ja5hQ4w27/DfsWD88IygMfHKs3d1G+DqrJLzi7WF2/d/qFfDyrLP8Z+
tqMgk7K1+K1bMkPyNjhVOBrwWo2UiWOpB2B6EMhV7S/iaM3OdpoN9BiGAbgj8aNHInx2Dt9h+dgL
39uKC9lz5f0Dkd+R6Bm9BktvMB82HjgivSLA3Theqr0Q+lq5JDLlr9XfNnRdLaEfqZJVSPmE1gTX
AcRhJ6r3VFcBj3CJv1UVebfBE+DnS3daEpl+OyV8shJUQAjXPfzu4u6Bc/rvo17XuQKa0+Btt1XB
hF5Y5lZsSNaifbYYlR1bRsUaD+OBbmGLb71QJiFLrluaIOa+0Z0YvHtHYk7q1eGZVHqjCH/sbQWV
u6P4fzxTqV1qoQbWgIEuDookVFzJx0ktCOun8kljUMgczW1RaZZX7YPFCJBm3V6ihGfFy3xOeQSU
0fsTfCkzdZ342yuJXe7q92VcoC+D01Lz1FGRyBbPIU1i4YaLs/UNqFXVIlFe2T/6BMKQfXbCJriZ
OfMs0JQPwW6zMjgWUhrippMkXZYP1XZ2a2WNAz+ojh94ZKmpUCt5NNpgdNW1IGXFkAUsBJCWkaCH
8UktXi+c1VDw9zoFjoxVupaP8FsCFfWljAmWRL0oEjOITA9+gEmIbraR2cZcatBeEvwtj69LU4By
e8wcjhkHqUxPr2GVnQXZodCPIaWMz73ahF09Vu67DXqJczVJCMxQY7mfxHMUZkC7cdhKtvumXe54
U7iL8xo4gkBhtV51MgtPzw4ovt1reIwJDug+4fUsaI7PAKDGi8+Qb8npnjcJ7NEi25Y8Llzfbtzb
rOxGF21rS5VbKhoNn4Qoemgn2JBYG+D/eMZS62z1dKYvROWgrbSSUKL6JKzNGhQucy44k3i98bfC
vJBY20e/5zqu8bZEsQwG+tCUfMUEUggJnLd9OUpaAN/lIiiVfoXncT1NbjEWM//x7kcC3CdpkxBd
BuM8M1JxIwrpflNtCG/SzjxYABcqW2P4K7bSiF9TZ48XGTPf/9+2ucmfMoJAM3j3uDGLFadF/ydk
R3doHvcyXRY4R/PlSDwjIjnZG6sfFm5lf02hHuupEaVjA9AvvskoO+6nb4CQUYmlXEbDAW8E4K/2
uf8KzCeaxuMY2knm7q81Cr/0WWhyXRnX2Kd32PUf6GRvc+Z6xtb5HMbzodSkbQHLRGFztVI8ckg9
kmuuCBHw1oStkq/0IhFKSjeJkgSqYbCgL+Ytj/CfADjnH2wZUbFcZGbcfSgZzS7t8sz9YFcfAVxC
ArNgWzGVNbm7dqrNgtQBukjAIu/0VZJdA8KRBOWZCd8Obk7rf+VbB2J0OA7yr7V0DjcfC30/BWQK
GzQZj+LPEABfTHH+ySH1+xr/+OJw+vK4ma6sZg9QzkFjSlDSc40aRMaXPxo4Iop+qBiJqXuOgB1B
OANtODdSeU2rQjCqS3B4jjI9lIZJWncHjL+ulQeIOUrLW6cxgf8G6D2w+yoBzgnjGFw9l9kpbJYF
MqqPZP+X7OZz0Tc30688JPvFaaB2EVGWkOISB14kw10Gdd0Q5RoH3DydWBNx7KTKWHIeyyzmFFHJ
NhU5iVuZFkcbpcPVx86LKreGyokGQ7exDeygchn8NGnmIDSK5UDftIzYYdKBEMErhXpP9cIdZUSt
9CJmhBzIhsRs09QD0DIXys/50/nP0o3cCXCDkBBvyXUtS+ftWTnWMAaCK80mI93ek82UqbFYwhlx
yM+lJRcdUgMKneusp8nUyJIGDLjMFBKei1h7FMP6uYn2bxMTuKPc31hh4HUi6nRW3nckPHhoVoCb
R/u5TzJKIFM3P2eoKYQyNNKsvm+vhfKfbc5rl3k+zWHv7OzUL5Vj7GgfCdQJulYaAgy3sOahiauA
41QtX+s8J2HssL30tS0dLScl0/hWBFsQWVdooTOgu7T0xRK2ZmTrQ98sTYHkX3NSmTNxiFwbd/Zr
/blMEM2MMaNjPvU1jmccO0G1/mWaNc9Je8AiSs8ik1M6kr3quZaJKsbKLHFOEsP+VWqWnevn8ufo
bjT2a+k+MP+M5iHvexD8oH2W1yN3tAC7ztD48L1cEEkhHJmsq4dJHB8/FrvCrhSWeXvANSF8DLBk
KgI8fWPcpGRxtLZJoGCdaW7orGB5yIt/BZwgoZdR98YEkIwvP4JCOw4QgCEkyaD6d5XWBg942mxs
upGyu/Sg1ev85wcxWIcgbfAmu5MZtrNbQkw3VVrRs+0vSkbaG5k/A+rMQLP9k0/7pVj5UWj5wQoI
Wgu4Xrr/GPd4LcG2Z9/sJD1fbwJgw6q12TAUF0xGmNf+gENFWBATb1wv5EJwF6su25YQuUQgBPui
TMyCcE1irq1vpj17RSW+jH7/AUCmeX5oafF/NSSC32jmyMpMCEhUk3dO5c8rCfE2nddx2d6tbjRA
Lo/4rqbiOxfzHLwExHFT5gfCEP8ED4gbBdroJz9OSrxkALkxlsX2vu25adCjlQCvB7zSYXTtnbKd
ns0FKHvUsnv6hcWcPNGHfH0OhWXzP5Pwzk9aaouPzRgikiP54+0EQQbHYoCG7IYaVGzbtmo1QkZd
wEdVG1QZQUzN9Y2Ze+3a1E7THDDGW0QZEBairrnjOGpaJnvEgVhVygmnn++sYLwVBdO8q23WtNhk
RO8rYaVgPy9eUaCdwG1I98C7V9QfGrekLsmFPd8swaP5ktJU2YoHYh3UJIbRFrsy+wGRn9zLvq0N
O6ME+SjeGQX61DoYhDhCxwaKxAmWMmlGhS7xvZclq9rKrlxsRaMa2fJIEuhQ6qAlyIRM3IBYfGkA
/iw2nHjotCncDed2vomr5VIZPlVoHUbBrG+00R+NYztIOK6z8y1ztoa/RyCAQHK/V14WnrjfLoN+
pOdgcnTzeWAuARsPH/c8Bk3CGzv3JcNbywFX9DuuKpF1XqWX+Zpe0VrivLI3q7lV5HanjduXe0+F
bO4yNbLg5dIFMeQNnu6KuuCrbrSAt1Ncg7/4z8PIGg7M+A8OIKDMB2k7J7hEoL9MQdSPEf4Y/Rg5
Lbrz937sM3ayOK6RwRNZK6Ep9yFE1VfAThbDZWec7Xtb2dCEvJ7/dnPX8QqHVHLw0EMY512wv7rs
onxDvkb1RYLrP2DcBJ0N3w1O/pW6HsNi6XbYSHLdl8XIa2Pj83GUwjFutyl7mDZVHmRO5m1n4IQX
2qB58cS3g6fG+0DoKhLl+xHH0rLMedI57Fo0ZxMaAaYmLgNygSsgI43QS8Q1G1KGU/qGcuHvcILf
8LImQ+UVe8bzBZFixmMLrr+GcR8q3ifT+h0+pP3dj3MEyKcrrKmJiR3fYyFY3fLkmWTcVP3Htyd/
w0Ov72eJwV3QyivPxAq3mW+W91GI6KCnNibPlZRRM4W/p78KQHYicUalzwP422cZYLlGVcMbu+zm
oTUXMqQJlUY85hxNMlyK7TuUZN0B+bb8DImUINCYQzhGKvsUFz/ISoMkIOpHzEr4nh43aBQP1Mmf
NI6AP6QgEa9j0EveTSlqEkcONkfoc3JhJr13RijK1gn5TibM3YrgEf7qjgG9st5gGo7YfFrQ5uH0
SvwHxG9hNpCvqxwfMa1T4LIn2Jt5IUPAKtq+LziSrVQuBTG7j/3cefRb9bQD9YYSu2f9qjAzTmZS
PdjJCK4HI+xpa/ccDHB5gsljVG3sDUDE2tth+FyO5FzChmjJXjLJi5aFCHmjMW0peKRoFSD1Aso+
Qs34L/HOE/JyJi1G3+p2Tb6HRm0Ulkzzfrdk9aM/s3Nxn4aGRhWegx/+I/zT8z66fsyg4NesM43H
OyCOQX1VOutzHTYbkq7lWOx3oUXiAkQsrbsEBZUui/+B4MaXeBLE6Qe36T45P2ePC+LY2gqbOZds
J6YpB3GDs+bo3JYPnXVnAzGys5eh2XUoRTafsiPPIJCsMnT9Ng5RW/1xj2+2xjHRWYjSFnNJPcmj
b3gXNgWXu2WJnLFTMYGv5f6y1P8JBMuYi2rmnwPTuT/loHYnSFvZAnQRFrlC1fUVX4h/pmqr94wi
hX1ixr4qiuM7TIGH/Cn0IMuPugZwofP+4r2qbEOiUaryE1QQxFnrlUAR4Mx3qMqhXW24RaGKh7NP
SqivnpYEfZ+dxiovk2w9jd0LSmptZWCHS6IyHqCpkNJ/Lzu5iYLpVFFqXgjPehYiiOhhrA3gUQcw
C6g8fVOIZxb8g5Ouvlk4BbM6vCuXbGeCm2AJL4bg+B7BzBWLCOUVi84/04ZY1lT5veAjiMs5gQTS
kfdAnHIvjEmYQjjrF7qLZ08tevx4Mivn9+VKUcT/RN4RqMBKqfYfmclBV+DCMrZTCh6iKvTD5ye3
n6DU5MbInmVKAIBOVlNOixRwgrF/GDsfa/XAvB51/ROVKlQky78DSdPwUA2kcucwHpJYBb0B7kG3
8AYQqalsERRx5MuRW7SK9ij8eF4L3VmhkLZQkoCbRvjzFXBc22FgJXQJa0ErKN2q0kRvh8zbl0Y+
thrmvT7vENG5bPa8SH8L/6MTC4/f4YmR5ZHdqMmtGYJEkGy/xuMo8SE0UIDwhxXdR5rD/JUtw13S
ezcRP3WMWIJk501sqWkYqsSl+d9W0mMOiz0dA3EmO3+Mt/afYin+bsKACpckZh4/LzRcuhSfNLui
IkEuboBuD04kshIVduHgi0d9tavOuJ2Edqr/Nhga0ClucnN0LbskyBmS0+k0VYL1Ik7B1veY5BPw
Uu6y7n2NSbon0GTDuXWBy1CPsTBDxDZoMPQW+ty/CblKzyuLEDpnXiQFENhaNy7HIfXNC07K3Vk0
JDkBgt1pC5da36Xum56ZEssTiIvSCtVePgebLkukuZo0/6/oQmD93S2ddJGy6Mi3qQjUSoxisnyI
tJBpiJpZdmXcSCJbZOSDS586UPRw1yKiuvHNlVtjwQtXtTYB5ov19s2RiZR6jimE8ilXxPUQHWn3
9rxHQkf+noDDWJedsFgOIqSskBenjzslVwQDcNivkpd8FZShK7Mw9FxhS6fpxWztu6l5WBeXrubI
MJRXpha3gwLPoNb4NOZVWY+PqKzymNqqb920FHA9LCK+KQrIVzDanBqrpOpoiaDYHGuOzcC2PVPS
zCB8BBoxhtp1/VdnJDH28r1rl9i348gghwTT3o35rFquhhgKEvQjQtnYY0bCaJTB06xegfSvGFv3
KOY932kmilL32X6Rt0xumrVr4pgp4s0CoSbVaTz+3H7/DZSklx6I5rqscHO08CySAEVXY5IrfoDg
JnhWi4myDKHGtBl5mOAVVWpLMJdL2aKucD1gC7S1JAvwsvIBnUExsyMNmymSquVDjr34dLnNbs+D
z3Q3z6wPNyUuIqGB7H7doD93Ghd+PRfnlxX4UqUs3X2gxMcc5BbQWITevg6JxyV0u3FTj/mKL25B
imNDgI4ul6nop47L6qwTyvuhUMR6LUFErCvwonI6WCvrGGuWkLm9Z/v48zN5k4WKC7ty9/vjpWkF
SVJMsJfkNfXuipyYkKvVdizt3geDtvAT0mUszwXQQFvQ9e6FAJeVLEPABzrsgUBPx9wIm9MvP4D8
sZLaR9OPq8AA8lHq3K/3tqgE/4ZqqX+hnq5hJVR1q7NqLOFLebTinRY3nt8eGm03pDzhcIKWiQ30
J44JKQ2UBsgGRfKcGp4CglLIwSGjhSevELPYWnwsZdFxOf03LRHe522CM+YxR3iBYw0X7iTg6LyH
+IIBVmQLR8hpnaRimYIcTIZ7EIVwuJSNcsbzWiFWRBw9PZBOrUPPg+cqLACDOFrP4k22ASadgycB
lJYGZ4AdcEtA0mf3foAoM0O3vZVikAxggJ72j6L/7AjvI0vHV+2c3nWj0E7WC9fi+0wRHXH2YQ/L
qN8zUHqHkfvIevgDXVv8W5vHlWWsbkHRisW1O/rZ5tos6txaed2bItHC6H2gsDZzGy3aLU0o693h
qLxM4PruKOpn37an2GSMhiMDn/pRwh/wqg3GNLyKtwsPLdVrfAZFZR6TZnZHVCsXTVO34cojR9C1
8mLJ8rKOLKFFTsOdQHAzLas8JzPtfVWO+sjH8KdkgjdkUUBJTrydP/kWjGnAKdyYLbYMYri0a5oF
59asTe2NArpGF9YS7X5aAG0KUnYZeo4L+vWHg04INuu27Hyb8SLuONyrMOxWV1zRPg/Hrga/w6rx
Qji94lHy/L5Fb4TmB29z/0UlD63v4zoOGh/XVlQ6dbnED4U/t6AYdra3ccJP03tlK+hr7fo+ThV4
K67ksAKvJKbhd6YuJymaAB1eU0IlgxceWElVri/bWa+GCtiebbDKhX39KFVHaFpF1vu409hYYVYr
7o2KkZUYzgFLbXSmVic5cbHhm5KdQZSdeOXH7+c4BX6fZY6nlM+V3oUMgUwaHv/Aa9OHeOVIYcdp
W09xDbabylLvapRpkonE3ju8YUo82NAfoVe3MDN/uXRRPTNo7dOuAtlvOnwjDHJVug7pW9v1+qIm
lskVl48Kh9i3P4JlheWbySkDkohBv4TZnGyGnQi2GFWZnoMDGm4tu/4DCPcVQdQxg4N6JU/2OvfU
SSzweVW3o4TMOum1jyetUdSCam+tNSX0EQ2WOQbyHuKjjkJ9bnS42sLeU7QHj6X7Dho9GA3gfYji
+SWbd3rBZCy5OzmnNbPrBWz/HrMqq2E/K8xVoRyTTHiiSw2grD48m+DzZE64FlCEQommUYqc8chI
McoyOpja2x0ApUDWWQ9oN/Ht2GqQ9N/UtwxOOxdtiBRb3rbCpzSgTJqdP/YIGYrnvZmjeea9RjCo
0WUCdJ9372DqLTAtjsiNTjDu32YHjTIPdsbJ6Dzlv35sQ1lfEGs3trz35gbDXxxHkIzgpTO0oaD0
aa7jUM/qFhy6MEL8bjDMa1ued8cUtDTPpkxBQs06BmklghkB4Q/+5koqdZmSQv/Cc037bO/XyBTL
tKyb3GFyrxgiIiXQwJ81yTaoShdQp51Xhv+1MXpueCEUOfYs+NcbPXt/KQ0FJo17H8nKvoF+jDxw
ddDamvlHwwy19UugA21A8tOoxuXfz7UyNGlYCI54eOfetILmoamAFxpmSmuUTJy832bBO71YGT7G
2Q2/2VOwG1lKXpCuGOpJVMRyvKx8V62Ytp9cljwgcAGA2/qqclSzaI9Ybm6P/0VG2kWJr0jeVRUk
KF1i8v88AOlDtXB+F+c7XVs2D1Zf0t+5d9upKMvJPFO7E03VZpYH7agHQyi7MrfI/KUONxN6vnxA
oqnhCiwtxq24xKygM6rT2gacDp8S1AwMcciFHCVT79c8bzpRB3VqrT/sUgjXJFqZtOTAq5OTATtI
VoHEcLZEBdCYo9rqAwob3Nd+5pQ/G8hW6mOPsGaTd0BkWDRi8QP/j20SJdtD/al7AQrsekJwIt/9
DOxYfWGLxzC/JltOK8TzHv6Qcgk11zb5c89jTN5wtmRHEEHHx2JI8Oo7cJTSPnm5SrXjmtcpo9sG
FqO8v5dNMyuieTNN/J7ov50pgNg55Kv71U1Zmbbwh/frpFiUnSDPsai5QeIL2V45coRMrnYHIW1j
stki7ishU0IK0bNaNYiifEdS9GNxiQhKfuOHtlFvEcOwRJ4vRHavQ3/fmGjfJqQ34mkvAL6zRy3S
+nJypqUqTA5ymZQVi2Lh+VdAIqJso95COwtLRBakSWxZAPPKL6RgQvIHERSuK/gvdkA0wfDnLs5x
ZRNPMfLOS3YZwUJ2pLuSjkCiO74sWpOZA8HTZar2pbjZ4smCvHdKIKl7jYGIlfwhqXhuNtfkcobJ
35O4xUW2j8aULfnMrgQ2GqUpJIaMeJCXJr37UfbuqlzKd5YdkNa8d+fN8xzDfX3aDPUiLFJC5J5C
wKozpHw5qt0tyo66hV10cFmrG8YK07bG74fY1Pvkyop65zL2Bmpo2QnecsjZwxx6REabdJIx+7ND
0FmQFKySIe9pp87CX9RT79nfOBWeA26kxK9uLuDz6MDFq23vNpFYYNmjuER2T3A/W5uFzqmNXEqV
ET47ottE18ORv8ujyoufpq6upJYJsG36WHO5n+o4PzlSaQUXHaVEBUZzgcRdk6bU6P2oB6cgXB6G
3GyHVNn3xS/JeRFjNHzz9FrkJlGFOTMXGWsdTWQ3FqXF8LRFLi3TXImRdE4PlJTW2eBSh/9rKLK9
0yKReKwUo7FzxLI6Z1e3bp808PmZ/LS3PKjOjI8hQZiKgvIHdTcZ62wmlP9co8mhxHXHoxIUrESu
FBA43Ab5U/QKxXME6oDAS2IXp7V8MDj/aLDuG+MuwXWEEIVBhfeRFFoGCbE2HkFkJfNSXN2TreTw
ZIxGa4/GKhtTTUTnTnGelLpR52GCdsw05Z/OKiEo9WaKu0B/oxJknAkue3g+YO0p+1JHUdudmGZP
7LwPRIaCwGO3R9h0PJrf+IKv+RY9YrgTgYZrAQqVUbimuJzOCzUBCbVZm9+cXpnvg/j6JUklfysI
hc+cFuRkmJ5nll0wHihhUaU38nO+JxVcMhduBmY7uWfn0EpY+yUqddSReRI9qOOF6XPRT2HXzhk7
mIEn8x8VDbQAy3c9b7kNkUHPbfHFQgcFxfi3eFLZbVX3gyeJO6m6WnNxNM6uSFgz112M9Mtwbag9
xxN6rdtvIkCyr7Ybr8MUImYAdoQiDUL81qQLhoSKKlIa0uwfLac9Eg1jb0tXstmmNx4UvdnhJEnV
1751kGnqOC8LQPfQ1jPbiFv7Rm26ht9LqAoiP1wHI249fvp8lTT1RQeEy3P614ZkIPMl1Vfh7Bnf
kV6SxiB37cYCo6JGIKn4XLh/Q3xwbbUDTj8MbxkLde9HLCxiVPnFhXrhjaYrvlHMEIpkR3Ng7DXA
l2hbl/ShNMFcmaQGrw/+HJlRS6zUU5rHDjqciixakyJlOKA4tKyRVu0kMGBpByfDXsEUL16Ammgl
1t7k0LxzOxWehpUuBotkm8rGDUVX/Lk3CmTYmByeX1R9SdKiFJ7Tecn/SF7+N1X2fv33E65UdE7t
iAsbLzK0hJXMXPzWYL7ccJ+pSz8XeQEUJ3ue0pVa54WLGk1eUjWCG2/FBjjIVkxeNU4r4SEHkCxg
u9jAkyR1Seg1X6sYCuUlVGHTmxYabwLj6roL53+5EzGIf+dblwWjVVpizimSzy8bPLYa7YI4b5SU
eSE/BqH5gyjQ0q0tDYhM9cvLRlBCd08h39PdCGTdIteVLPuU5YTcxTfdQ/PDAH2th3bvAM+BhXBA
N9PUoTDgbB6zvDJsFawMO3D61m9XwFOcRiSnaNliOJfea4NH6PBTviz7iU3zLQ/opSq/etvi9pRY
m4y5La2W6ba5zeHBuNTs9GWIIM+mbsN01GnVkXoZa6SQz/pD2K7KDxyZZVCnMhSPBBIQpSMuo3Gm
SDK313Kg43Jf0yDTV136WuwRGmghT4PyCd2E7WgzwsXzP1f8l6aJM6dRe2d68FFtG/Ez5gFe5nIM
rTU5/IU9r86YIAIOKf0BFQfKC6F4t3uPKQIoHgfstIcOjkdZEea2+534SZetkVwJooYfLdmVxGJf
6LMirDvZufaFffs3dSAVnupeBLQvQXnOO5ZSM4uakDDDOo3Pg7H3FWDodfJa2l/RFFO4vTqnwl3w
KuForwT4TxB9dluBhiDFkXJtLAR1qbzoVxNh6AzNaPRd+698WlM0mtxlgYCCs+nE54p7KVu9quy2
qoWy2zq+KtTdFdQoFk/+X9rIR57s58hzQuj6RSNJGgW5HUpnCBVygWXf2oM8OPZvMIg+KJnycsvO
sr6kZV0SKYm4vTr0SXEeelboLvN/KuXerHJaTg310DJcXXHfQr/bqs7XvTrTQeC7CsBMMNFRr6KD
euj55XmSmQcCwKR2WyMgq1OKOtQwec6czxsQMxUz2Tw0kSiIPiXZOdJZuA47NLX+UIYyZ6TwbTVO
Nl5L5I9RoPSlkmeJx0+rVv8cqISc1BY6iBVkQapYYkW4FJxgqL68dCrfgvHTkkNBbTEJGT2ijgdV
rOd5NTt9kzCbZKwWo+zT1BcVySV0z3GQ/BJX9GiFRgO5F4hPgLPknu0jun52KiU+qbhdWzlCTtj/
jhgbG3PES4ceaAYM1YcC2b2MObq87LIL+c8HTV65Wc0Qla+o/6xJ+mhxKvKqQ01rwiii9c0WCEBL
J3kBqWUG3Ri6Q4X8idOhCUle+2acwRzVbtVlxnsX6XyUT+I5VzMivTSDDo0DYtTc3prwXKaYYmGp
QT414h8jh3ChF1mXL8ow5aQHca/Gbmwh5I09bYs+TOu6Th+B/UXBHzclZQxjW3mlNUCh9Im7+snX
nSDnKMU6f+7BoCBGf7/TqMne5WBKRU31yPXTchoNBc8jWrFDujArATZ0R0SO4vO56tCwf/ozu997
iC7HOSWxsKNPfQ0E2AuFkAsS1mtwCykTHQ10RAVRnVKugDQ75aVVbkOkHyF7DlBt/46u8Bt10cGi
aQ6sBBuJZS9ywTldu7r6Lh34fKeh+yEdgEZJp2Yn9bufEN+iMMYyyUv4fFfCIf+DdjaTKVEvd0i5
erc1uy6C2BFSP8CUZcjtPO76dLMYaKT9vuhckyAfA2KPCdkMZVSjKc+IvSnePn3BpBwNrm5ctBQ6
uvvGzcArmpqJYmWG1sZmeQ1qPYH6r9BW+kZ7FRTymfm19lDP110AAzbbFuJ8f7ZDENHmOiJ5pxt2
BwZNAKK1Pm0t9xltoLDqW+XaIrmvg/rFoF9ldZMc2lEOB95uMSzQPy9E4PTHHkLxWTK63w5k+y+c
lJuZ6diAoFVg/4/WUbLsf0eHPCf3oqfvdGVVG0C9DxerwySf2MprO0Hft/spQ1aa5mwoPiYbDo41
cO5zytkQzMgoFjA79dbdIkWr9ajzjqpI5whBtvb78C1FMjjz79wrUwCbZNYpXj4tcAuqXYaih3nB
raiWPElhwzgfmAP7YGTqQO3x+/KCVBeuJLOo+BmBPTOCiPuotxCYqvDnAu3jWhwrwqV5+5kqIZBa
3rSsQ8Arpw8RGww4aVrcXie5ol/F0LNwt2IqUS/ynbxTeW6EOfJ0JTws7UNcDCtub3RjAX+2g4zk
QaKDJZ8MAv982KIZG0p0lPKDCy59eTMMLgbUZufxrO4Lp1LJdVMT2iWEQdR5alZQJQ+NC0JjRxvP
NOibWq/8o2n4mN+DLnZ6Z8BWfsoeLHSSUNg1u/6plkH9woPkkbL61bqRcqUlp1d3mwZ9e4A2KO1s
kubpIYYJKSOjfI7SVYl+gwkvGD8/heegvwEWuFIWq8VRCrY9BL4zzIarHfCZCtYU0aEmFsl5W5qX
IamwkU4wITFzBcKGNpNJHJN51mEST0V4Mr38P/oYqBC/DwTeVefDbWRRFxQIkMzJ9jlDMSYKnPAS
rlky3HXoYfcXW88sjxuuRkaJ7UeG0RJy4JY6TB5beTTXuTHd39QfNHztDhrYSDdT4i1ACKzAk7EZ
GxkvriAOLDyPLuhkXUceXKeW9sLo7Xksot1c1Za6yO+5feJkM7byZ3nux4EDgwS/3SgOyOIt3v8p
6jx2vDOtE2KMSw0/iHH3wUuO0locxsXWhC36WzMWUjlSb8eAEaK3W3BNsJxqtJe/cJdeb9GsLReH
gOV5AMZusCgKfGugAf/VAKNR1RtQC6/lS2ri0YENUZOL57xFnuXr1yNBaz8nqOJ0YUdigDr77PLW
wtDURP0NCep33uYL+ro+fS2siT5ND/qWodyGmW4epEULKmB98qmCY2Q4TANLPhz9opLAHINT1nSH
qVi5Wbw5U6uLeycTHa93fXn7lb3j7KtHq0NNYc8mgmBN0AXlBqku/1DZJwdBkKtg9g14orG8vr9g
nqcjxkUBZ+4turjDbKgHSOzi0Un8eb9UReYUvc/vmBXfy++eegqZKfmDYoMMcf0OAV17KNWQbI0c
G0/YlmHPO0udHDdt+RP26Z1jVPM1AgOp6OdyY9ckAHJNnq3cCS5TrfBgDmSVEDeQINfGbQJ0LdXx
3fODFHcLg9VKURkBN12LfHgWBKlXMLO+DJXoBkYaNFWLT+aeLdP5MAlOFz6qQCkbRoMTSEqhGFyw
Ms71H3bU6xyH+Ru9mIKQ+8nG1NkIiOxur4gy7g6GKrKwQvPLAD30ZaRFra11ral2g8FTsydXonca
AMVgzPiysz2cvr7P0wI00Brex8FtbTOZbIldyr9AArFdmTOxm4/CzYgiE3yRxJcCOd4Qyae3nZfq
rahVWrxBPZDBHCCkM5XhuFFj0tklFt1u8s6sWLs6Q+yUfzCQTwUD71ZLXkAVO6F+NnvDAufBX2n6
RzJMvtA+PFrKLTuhMwaIc2LNXQSeaKPyf3R3f3AFJoVQdltUf+CL8AeuUxEVcpi6cjAdsgxcIQ84
HMPL/FOteH2HwcqhePHQTA3kgN9OMwPAv9a8yLdI+lodykZbb0jY9jliF+eNnZ+Y1dqlblQSlDgK
mb6eUq984/OEIZCQVjyf4pB3d2MJfers4lPzPsXlNdxB9lHbj48P4FwTYqdVZNnhzEq9LzZQLHiR
D8EW0I5BfmBHp4RDnJ6nm8EL1I8wv37sjGjqjrDKsehqH8hA4SPypgDYhAlg5BXLbu4FtOO0pvSb
jtYh8p4Sx1UKhVf8ozAJnMRTKcvUdGfWyTJbfQEwGxm+TO+rgYb69VxQPNMlccGRwTULz46yQhwY
Bza16nCQj4fGCljZ2jklEjabmiwWj2S0zLuSysdr7MJfvbqVYQm+Rqbxed/yGvJRigyXoOFcEZBg
DiN0kuTwhnUctk8ChWVhdn3VphQAKks+sfglosg61++lsS1ZSpxsu+03XGiamsw2C61s+Giv/pNp
N+YiULt5U/H0pUwsCyi4nv069hQqpezt5cx46Mx49a0K/eB+ueSmSoh1ccZKBdoYxIhoR2CNISYr
5HwRsclglsL5OwqpbenKCDHDt2/jq1hBLpDwBXUjnNZAKFr3+rWBmNq8uff02l46JThAGSOBQRzf
98uQ8lZteHBPy1hqMa5z9ioGBd3mPfEOEQimRA3V+oaFcwQMWEiK/g0PP12hh3lrpcrGUYcZlNVN
kUYO6+w/0dw/bXMGkd1APeCCQyP+xhE8bjqDGoEE03jh0oT29qquFUFCrZWJIl6sXDqfnTS+q2i+
pH21QSHyEtcipsTODXCmymVPaHPF/ycD0GgftgFeSTeF1IB3yQRnJNEJ3JuXwDORpFokjuy8GwWU
DImU2qlHQNE6Bya/cgETMdYAlYf7VgFXgPmku7aMzNKgtjNf4jdXHt5+X84a/3MstChO01V3zVxl
WzG6ijMPBDF2LuOax3WjLvYLnx9Hp9R8jGCkUEZRO23pGQZ5kEj5EOSWSvu4IjQU0hdipiHyPc88
WrzHUEtKS5L2fAnk1NlNARu503b8j0Gf6pcAC/jwY0D2BBanLhKkLeeA/t/4z1RQJA+oAsf+nm7f
0SA1UrJ/PIOJNjbGzDERATvzig6agIPPKrYcTkxHGYhRiwQg49qI0H2D7M6K8gykdBHUzZwSRI1c
hFGE6AM0Gvhh8oiXbbybB3W/1daYEDHAbROknpcUDosP9Y1oTf08M0i+aJ/2wJoXY2qP30WgFD/X
MIOUAiPzl8hfFTiHyOtPJhFsN73O2tSd8bVf31kYrO3qMXcd8K/JmRCncNxE2P8dA7/JhWKv/Aeq
hF46aFfGJw5SBz1HiaQ0XZWetQUZ0RMsguHM6QHZBEU4sNIPGfG8A97Hgg5SAa7/emWSK75nyWtx
aTKkPqKjGAExLVlubf38viyv0taYbaNtf/BBB1PdU0vFnv74L4AW1FLF4GBihKtWg+PYcByWqzOv
lp6SKvnNoUx1nI5D45pbQ6F2AGEnR4ps0L1YfJeL2ou2hp2Vlt5CmbRiReUdFxVDbi7uZI1Dbh/w
gKcx7pi5BNIGQMoZGo5h/u3kBzkPCFOrQ5bM1R1Fyf3ItPvwmSj99Wv2NsCgzrZ9V4/H4H+Mg/8a
eDVNkLIOE0jiDjM+ll4Pv8CT5+e4lf5/feArhve/yV8YpLYcqRbmT5kFCK6vWRDpGS4BOzgNF2XE
9wcxAmgImAu7kBpH49eNIlPi/xGCbHKsCGx2/px+zM76gt1J2/W6phfpYTvucRFZnZl3JlhaSJH6
nqzSUjVhbahp1jTmAwIneZBmyX1IQtg+NfOzQyC79e+PFAVGR8sJRCqbzOSbz92PkFAEpHp3vbJz
hHqK3CrgS5wPVjenaHCil7eZPeL7MiQiIWMbZdrk+h145wR1r1WxhPIv2X82/SvT2rqGEoLYCiub
7RzAjC2sJ4i4QPeOzWta+YVuz777BxzQAuUSPnyEMZHoDdmAERVkd7d/FDrshoSTckTjpKn3onpB
hn+YOGE5Jk8fOFUjvQbRqa2REPdl2x8+dqj16QNQs4DIquQW+plSZWs4qltO97nYbuyYyUx3BS7Z
OlyvEeIT6c+L/GJJcYogqiIBWtlpS7/85N+WZZUmb3J+S7783CC9ctmNaGlXJET2V/JjTRwn9vpt
bIXrTaDAabD411C7wXAwcdGZYcYDVFuWDOj11VLd+bRXXfp5cO/R5LOVsM/ptEBxSiSCjx65jYU/
5cjCSolFTadbtfh3T/rwoG0gfU6gAEYZpQxwWMXXAaTnFhAULwpYUe5OmLjciBwzezYn8XZQdEZj
VN+HhsTbdmqQiEp1ll/3jLjyboZGgZgLZI7AdgZqgnSswYiz3MzdBb/lIpqTgqgRANfsUoihegog
UdJwCag+VoZHZu3kJjut5ztMDWff6A9yCpREqJ8OL42WIoT9rviBu/Lms2D9Q0R1WKQX/WNK/tYZ
Awv53TCQbbY+CwyxPqp8hmzsDZo42YIS00jl5nbgIBTNGOmy3RCP/o9CGQoMY0uwOQvOVcrgyADO
3TaSZyW4YPFNCL+GJsF5rzvMzCATQ2OUvPzVMdjYF32YVHINV+Nm+7Yuhk7Cblizh7xRogitsg+m
OqIIupJ22eoQXmR1rdcGSWhmEoGpvU0eQPwGo3miWda428yNX1K4YDyqIpV2Hhd1IG/9LwVrZyvX
ExjrdlA0qqxnEcWSWhOX4UfI6gMmGwbcBvyzO3E7f6c0GtU1/kwY11CSws2xmttQsWVF1fQOj73W
MfzoOZ86tUq7mhGu99SkjF4Vtqejl1z/TvvmNI+7RZqIQSEWkn7CmqHFETlYFIQYtEdAKXl9U/xp
LXvZG3r7SW3aZnaaOMzoQXhQ4vvvzmzVfxzNwF83gFNEKg4bAQAa5X+psCM8m2YR36532D2hVBl9
y7fSZ9aAWV5DfjuVrmmWn/7b+pyXZyPKzWwssrScZtLbQdzwAJU8LbAujIcEPZ95KqHKY6pmnQ1d
wZVgS8p0/XM+c9Jbe9Z2hvCcN3OklpseTisMlDny4xAmCs/8fZNYJ56Q2gI7ybljU/VwBI7TUHl6
L8sMJ52XCLczlikhecyCahT+gSX9i1DSG290gyWnGf+qqvYTC4z7th60K/BmgPJEa8m//YDPhnR/
rCY5lUN4bHeyd8dMAHBiYCVvLRyIfd6ExaP5DPu2j4OPlHE9/ppHDt4V48WZQBm3ZymqUY1aDAJ3
Q6fZs7oX24KqLTmLLvH9aY52B7t6oUsDYPdeNxpamYj057nzjvIApPyEwsmnMoJfeecPQ8OYJXkP
yJ4Bf9VA0LdedJBtsyFx2rx6TQh5rXGt2kVmVvJfMNNRli08hB3ID4nva8gtqPPDOBEW+cMH8Ki0
FVnTZRi0FU5fgtSDd5+0AA5+w90OHth/ZuWheFeYNfnWtTpwzJTsMCTs3cSKodClIHs4hMzv95Oq
7K38lBsDIkCjZzFZ2W5sf0MDo07KeOZZwhvN8/E4eUWL7nn5UQo8rJXezKXOu8kyBjEJy6JiQDDh
ZCAa5nRQYWNg2A5nvI63gpchWyoxGkUv2lOVj5NmeuPElKnDDNy+snnCAYDzI7XejF7pHeKeDr6t
1bzM62ZU+jJ3aAjAsZf2rwFB6AR9OAzRPYugpQSdMAo095vSm+7R02NGHQKzwWSZZxcGFT2XqhF+
UmEIzTd7fVYUOmOinGlM8v6YbU/gWirnCrPAId8uXHKubqNxT2TAYEXAzKjOkyWHW8UwQks5MxuV
jUroqwdlQ6Cd+2uBVkTgMg3YuxhwSWxZBcOhQsWuFZ2T1jkZeVkT+trOjwFmW3MZS/QNhWT4kp5f
w7cpO0UIw0DmSNSty1fRllZE2fWjIhksbFmKnA3PlODN5/mbB55PNe60KqLH/uc3d8kuydrvFhB1
2tb9ZAHfQ83SNTn5WbiweDJXrau1SBkZ/D9hXHdWK/L2mVqxmTzljDRaNeEXWwCvxsO6SzcnWlmp
K3oAFqJCzMCWK1Io5PN9ub665KEhlS+sAIIXYqvn+gRCoGVGkObDP7LgyzhGQjfHCSa4M9BJO18X
gu+zOV5P9twNbWxNZ+o5Zmtj+GqO1c7ECHBd33DwHy6pEqrjHp2ABq97cRj3amU0sKgVek4z1mMa
lOKXtQetGZZkNXkUQAk4yQ28HP7Z0rOEAQEU9x1LiCFJg9lBkaXq1dRkzkiKWdLyKkyJIjY1j55x
9o8hgjp3zfVzq0QYt9JHXA6utoS0oB/tufsFpoFOCzrUWrlqsJT7m9C7r0lxipxmL6hDC9GGOwI5
xhNsvzFuaGAvnCzsmhVGpAjxkB6URVX+8A7Rl4ZP9sBPNKvbk52146az+ydd7ySOxhEnGLoI2fDF
LJ4Ah8fX+/YyVHU1wCiYsbDGcK0ZtgGRzewc4tY+/i6/v0ReyGxHLfDGebwLceT5zHeGkHpkMvuU
tiYBoFbx1KbXihG4o0E9fG3LN/KRuKttIgSIsU64KSZIa//T3yebFbadvF9Mg2u1aV3SHYnAkCeM
BpKb7geFXyL08zpvvMKpZCEcLy+cq7oEGfg7UqIPuGcRcnhkhwNVvM+KS4oszJNHfqoATXU7R20F
4t7NiHPW+3Nfxwx4bDymPFhD1tiad0B1/Om1YtMi5gtPnBGaa/+ZwuDH6l+HOTe1HVoxMPfoTNiN
OV94WCaWo9Q0jpn69wnSiUdTu40P7mDj0OW7m6cHHaXZKK4y/sPX3Bw2/sDPNehZnaIEA0ZgR4Yt
n3XbH1GLdR6QN9Qqd5sWT0DNk3IKIccXQfSGtYizyk/u9k70nrTlW4bKBjx6e75MQ4H8JGfDJzZd
g+dAEooDkiuWpozBu1yDmeDvlYmVtiR6yXZ+OfFEIYGmEbN1RAIK39dJhqK57UhEBtVWv2pECLr2
9SvC/EV3zTibh8qbmLHqD+b3cQVALnlSTQK+s/uy5o5sBOfozqYrsQRAcS7S4QznB6iVhHZefrLr
fGuZb9ekL8yzziffBuRogi/2oQqJFJlHIMSQbss48VLtBpHnSi/m6+aggNY4BHBH2XTr5iJNhCMQ
PJa32IbFn6ECcZ5H1lGDm6QegYPgZD+1HRMDyTccp6BuP/VRj2cjz1kud8NiAESvdkQ1Ll+ZZX2T
Z2ui3OnCUTWdMphgTPWT610qIvdTv2TadtlY2zCYfb8rFZnF4/8NHgXi8jQel8jymzVsiGqMSM41
EuQAvVpokMUZST9WzIxU6br2bBBeRodwx29rTW9v0+/vuyFwUbkOrKcmsD7nCkfiUpAwUgfSqdCE
IiJ5GE5w+EF58CaFgIVt3juocBAqfUlUTRDXuU0YfQeLnTp/E/tblBNO+7oWLWF/ftR9uF6cryM1
zcHRSSNu94+AoedbbcdxWAjG0GQqoVQc3GGqw/dFiDQVeB+vYIk2+EL8yqF9mpKZYVJYE5m82Kdr
bcWi0D7MbaYVzC6Hr4eXPAgkSpgTLwC6+BOava4eala3NiPqogYBx6kns6XAUooJqZaEHl7AneQA
LiKitcVDyAmbPlLImjBrBLVF0QwsvA9oGNSeaXRu2SAsr+ZBuZ57LOiqrL0DEzfLobvkyWF5wpRv
941Jd9+B1aCxOra0wxqRXUpfjQfRsv2jIzTjKMXQVua0z49ZMR9XzGgPMiAoGLS/2muWXIZUw6EM
DWRNjJEYKFQ0Jgv+mE2ZAQFzAFsgeWISFoUvAODd1Uo8m3KZ32OjMMvUbAiMVL9lKFbbGNYRmDdx
qmSgZhy9wltTeNAKVFgD8ICrRCc/1wA/M0Vh3FX5X9wvmOO1PQ9D2SDK/X7a3suX+Fo1zJiVhJMb
Kjmvn0ubSSMhl9msG45mQhI9X1I5Zm9l3tFR2nKFCrPaezJD1FL1LlA1viGJMeQPm4wfoj1/sG39
im9rO2zifxwCKl+qGtFIlZty9t6mPFFv5/yTdMF0Og041iCGA2bk/0chsDAPaGCTOXIrLQa8zcmw
aNDw9jxrD/m9xkaII8A6wa8zUDb28txqM0Zn+l/0OoDplxEAaC5wFhgVavzFX4AMHkTM+CQGnvgj
4oF45514b6yOG42RzmfCFtb5IOY2sQUd/9jMB0PrKAF7vSupzwk9d1tSKzS/6n6RHjNkkssvBwOW
x9swoBU+pKpJzw9NPjA8Njv6rTntPp0IVXufXKccJtp02ytirJHPAsI3P0mRpc2ckCMn9nZahYn5
PgkR+hVv56DewpxUe9w8OldhOKRZuZwJLP40uBz6Q67XS3gbz7+VmICgQr8zgI8/Lp9nagNuwVp4
vmZD7ZmC6IKSJRLbom4QVpuojKc8m9mdzaGHfl00opH2QtBep62dEu3AWRS8Zab7rZGR5Hmx8x4a
YXb3qPmuS5u4o7vB6tSESg+j+xGqM/TZxK5eMeaV+a57oCw2NsXCmgG1hQCxUFkYwcyRaGYZtbx7
VyPpCL6fDfHUnsbuEx4FkGs5aNJUjmqdyxIj3KcCinxvhMNkhEF7Fw3QxsD21klx00w80cFwywNl
zRtpGmKnLaSkofywYpwd2unn7pj9hrwtdHVEqOZVj5ROULyMuFpd9UC6zvNySGHfWdWh3/CBb48c
ZpMHkAXHEkS5SCKbMac4ovEcqgyKHTLqzsR0l4cB1OruRZc6phvcShDWfLhjXXcZSnGdTTuogidK
BJiRfAyfzQVBlhC4aTGFePTZnjj03AGHarS1aA3uUWoyhOI71U4X+d4eSrzaLsDEIsrzuk9yMTJ/
l9mRYsrirB+IIYP44nS8TDKyY0B37n3LcrRgX62lcW+EFoqhCoOoGhttGnZ6DyM3M+mXcFbnhXyV
kLyZC2aqmINqifCk+uPCEbDk6KEyu76YGxubKVlR/0aK/hM28znmgaN4/pv/dcWaYmQexQdY43P3
juZ9OP1d888bA11XJA2cwcfXZJsd//13RXEagDyzsg0+aP+JDdfJAfSSIwRDh+i4GWj2LRC2CQgP
qMflD+LqFjswaC7hWZ0DJAYfU3UT2oO+i9hb1L5HPXjQguc1PpQw09sjZCeuDb9ojZxSExya6gAk
fhR8PHez8O3zVwhfeur7R3QS+7CerOhusoXStF8V6A3Wq+aBnH7vRpYYWct9L0xfFDe8GeHCUZsD
ayH/PmkZXiSFaOfFw3t3NSdIeWlhDcGhgAkGnbw///bT2pHrCQkHr66hDU9ccXVa4e9WbX1k/lEF
3xmcCa8w1ArT4ZPJMEaLv9TX5oEKpUsduompmyNYTuhay16ZGdXaivKE7t21rL83Fm5bKVgBWBqk
zUsmsDnUj2HtTEkGyUol96dCNELNYfxXz4xxtAOTFkH8n3xd0bqpeVkiK1sObduJXzUehc04gmvc
vHvX1osc/ZiGrGtKMT6V/TsGZI6b2h7pC5nxvw0OCx7MDZaAndTGdHTmyDhn0JZbiO1iU7AkTBUA
tO5mphadNO8ZDSXXdG4LpqtN8X7DAWPr0ASddeZf0EUHzStOu2dklAuN215VtbCCISOuMUGKXlqL
jx8sYdoPOJK1kwWyZY5/CTq28r1t70p4kcuqme18xIKabiNbOTSkCMsceIcwwUuBavUcawrYut+8
nACJDqp2jGO3eTpBEdEZ2WxOPEbgKfIVCIs7twnra7CwX3idqCgsOpfkdSukMftMWiRdG46GR0Ab
mY1Z8hdunViJz4s1XKHY8G2IR4LVPK5K5i6vnrBJpte6GQuFfMAxn859PAyar5D9mIBF2Sk/DCEM
M9srs4nEL1Owc0+5nQzKlRDUsQzg5NgGVQ4JMlIy+hwSzzohC58IlRK6cjtfZhOg+7T6EZm700Qx
52zvfs3sJdjhMAfbiSkhFYl8u+9x60IFyP1EpirBPz/SHrD7tFoygs8g1rTWUvfhvncflZKsMjAp
cvVVspSGoiHM868izF5Ef/6ToeX2w00oZNVaMuwRL938ce9ppRXUHFmyGdImspilXS/IQMNctScx
uXyHy3X+eRdZutk9BDAeO165wdMxA93IlZoBWxjZLH74TDEKl7L4iDObwYWhUnxMizYkqMsnzVJb
3xkSwKcBB9RJ2c5dDNowNM2AbTRjsSDH3cfX30ajqdgYKD8rdsMpDLjMr/8J48Kk67br6vIVAIH0
sJyDg21j/FScf1hqlT6DFAfp1pydsnpZv0XpTtq7/UPHh6BYoyJnHB39sgvZIqc89nKozCNSTKnD
hVu4w6k2B/1VXshj12xQ7eKIbwdu2yofUlZJNr8BaWhzJ/jWXJNZCnq2dWVI6BqXzRXnCZt51HAt
zEg4+vo6FkW95hEpHapvgytYJkJ/hjC1RRtxBWsBcNG0SoU1cUP1dtpTI0pZwXhkQ0e0dl4DHfh5
mFdjoPj5fsCn5ZriVXVKM3FiY8Bj6CKS/NOHDFlFRrxzfemXBeo8J6uqJEyXlDudgtXjSXosTIrw
NzaXwSyUNnDIiKwlthnAugcggHCNyC77j6i96GOgV6kRRPMzrhgPBwzDkpcOkmyO578uShjFVqPB
51+GUfiSjjlYK6jRXCFnc5J7XELzTHAmF/So2hlNoiQmUCvJNzQktGvnfj/nTclTPqcXUPDuaf/G
MURF7Iq/4J2rqQGwL+EtbSOopP21Bqo5XNlLwgJsP4vj0s3HOWDebLxkL7OtLSnQvpdCRZJVZIs1
Ss51xblotMIyIdfArCX6QPQmXqOBtS51eLgHRXT33N4D6+kDQKfKqFS32FmXPeo7gAMmPf8wHGHI
qdcO4cwCuvZW/dGIVM0DGuMmtPD7J3CnHUcl8OY9kqQCTKiBMjMyTdyC3e4umBVIoZLr3wFT8EuJ
5v5vCU+9WjJ7J946/XXy390+QFgZ76T6D71o2XFPS2Qs9XbNrz+knQsicqba+T9wAldFoVb+dYVw
aQUc0FAkZNMnwOZRecAAUg++900nFDANMRkh5cS5nirP7L2whahX25eOJmE4QXLBsrzsfv+1dVsg
m/q4k6itsllUKYT7Qc07+J8ZmSqoe4JNWYHnKI6VKhe+9Xuo22t6v4NuoHBAKRrGFiomTP/CYDT9
IT/SkhXkkZhm5/iP6ZWINh2gpW66ooFtQKC6ggAwXWBtwI9djABxB82Rj8kPM6fjAgrV/HrR7cAQ
nhqEV6bfJUg+oglPvNxNFxQrLSp7cqChhUtkXaev0lu+ARjUFQp7QqArUPYMy2T/ixMslsNiRt0J
/L94fUL636ee+uY6urjFFE92vzGhr8E9iNQpF0L7NdcA95nUJQExRuId9EFZ+PniXWG2v49J7dNJ
J+LxwBuSv8D/hDcoCuqkVjLzPQJug/PcGBwE4SuYXHsE2auoWG7dv/AkMR8HHMPl8xLEmsraDysI
lQvSFwGb7P8wNdk6fxzWhoP4G6vjDOAqpFI6H5NOclXqylLggoB2qhUFwJ7DCtLI84c2fy4POFK0
S7lOxOtuKlTxraKgfglGnAmgREvHwTDJLvsO5XP4Yg17cIp9FZfan6yFaaUXS2hrhbvRQ+Alhq5o
YFRSXZ3sdzwiquS1j5Q85849gn/LEGbpkVulBoz9rAjRTKnpIKQqDbCNcUDAAELdxFCaLbtbKQWB
8YODOiQ4HjmtbWmwrRlKC98XliSlqp2dAy1TqaFpAANSnfgVNZ1mvonHw850ZJ7blMFYuuuJpgaG
hF2XGYVRzHiJaFy3fd7TbZSVz4NUwFsgVC0cEbFjwBFlxusvsQQAZxHcduvmqGwiDJxzXKZNWjgk
nW/8V12jOKdWkXvB6s9bQn5vTVg4YOXZytwPjLwI+QpBH3Uu0ut/wAzTtFSMjrbPzffxo3Dgqnla
jS/KzO1HB+ZJ6oUqsVIbATxrtgx9D2i05ki+FfUFtKZWT/Sjxd30YmPPHk2+aOV+2UvJpUFmxUYi
mkphoVZkkl9CgdEkevQqa2g4DD/B0YDkKGhWQp5cbL8Aisgrcr+DD1ugnPS0VnNt/v9KHKtWh+Uu
gK9tUT9qSH3+qiUbLdhw2yrp43UX3fh10sEiDs5EGYmChbqjwZ8fg9SHdaKC7LpfjsEbxp/5PkJa
uOsBMY/HnXxJ+XQ0ayClveuW6IUav8iAMBycJStd7KFGlXmQc9NQALbVbikuYG7bDgY3GZnGsk9h
r0V/G+XjaCM4zS4In1Ic8arC9k1OVaiI5VQJF8nKGKZkhRUPi14hz2QkCE03DWw9p3bCquZEvYtI
BrOeHd6kuWvKXOlsn8ke+j6rJwNJbJ7J1whP+dgkw6hQTBabFqNzniRvgdHJjhhwcuFia7AeFA0E
R8P8IHKXrrRjNAsE2iTO8ggEzZZ+LAWm2YWgWvCYjSveEBpaBakbt1IgSEr/1f6+Xt5I6Rtr/Cp5
xBx6OsWRjqo0x/0VQ56DROBLNIwGzBnTllS5cG6BDt19M3nB8j0IDCFm6FNUdUP/jMXKVwyuyoSP
ecunZWEPc76q/EjldsBiCOO39C2umqa9PmviL2j7dpytkHynmALm7QFP4cJsZ8ozaeb0MMVuStzD
DImdi1byjKt/UK8CD+Mg4eaBIx0m9//tSyJb7EyCUJSj55sPoosGDXAw45ol/WH8M+cFv6nXvCTt
OF8TqXKBvkfolMHJLiuX/pGrmuy2nEZnzz1howwvvkl+3PgNlAvjPK1r95l2NTFkxSaHYgYjYVRt
Kw5WO4HHPzqFhnouBC3ERUcDhrLRHVK3Py+zlTenjqX3z8sY4UjtPB4f4K3DYeGG+heLL5uUaym3
TbaBQuVxq/idNJvpVp0BYyr2cCzKSkWLMt31w10Xzb2mHlW76OSa+VGHP68lizBCW1nMIDQkrFp7
ZSgw+vOiC1/n2DhFGK2UDn8HLV8BR9v5idKrhCg9+WRC9zaZBR1Xf9KOxQ/8Pdr6HmCQt0Ryaq2f
+2fslegjeQ5JsMe/FiI3Ub/b8Bd1s6vajyiiK+npLNHzjHQJ1BjWmxHn5AVqQnxO0NNMHqqsQQ5I
FUsPEz2twh13d/mvLxLyObCF19OA2rNwPS0Wq16TbrOVy2kx0OG+kGaG2x8sWaClwwAMW46W8mot
7+xOEQqxhP5FY6gxo0L8LBrDKZFuRUfdxMLMBSr+H42I3WMFSw+CEKgUUGLP/y5oUZYhgnwSUSBm
h4+aYutDGFl0YqYzC3sMcS1ADRXbhf8j1cKP2adB9bVel23vs19RLfn4jM71tstzZFqmBXNMogGx
UZ4ZcSd+1CsQVPX7HooaaqRv7mkkRgtN0HjzpdttpckUPk+rA9fTxLrANqOg5gS+0s40sFkLbRow
lweelc9UCItVwqfocYy6qcoy8slLsWhA8sO7k1VaRbhpRVzq26AyWcSmm68lGBNavTLorJ9zs81h
tXCnDUDY02t0zwR7JptxJVwpeBK2QETI/vbCOrfx/dkXA2/oMBT/lyNeqfy9v3zvcf+24KMJiF5v
GeXIT6mOAAQxMP3OpEHQJQxTJKKwZttMgqeIPuccwWch2n0stqIoOu+QQ8hHXa4ZrUBnVLRbiomU
Y9D7mfovXsw72vlBcuQCbrrfZmyyBMAjZfwIP+1UcoZ+FRybBl7+X+k6a5hbe0Wz+4/xv8xM98ul
ORl/9B0OpXj9VJGmY2EgtvgeLetxiiKN+Gnt1Q9P6jEzdOC5QuNjLENADjaGL76EnXQatJwLShzO
GBJ4maEedL/XJT8nXHiZ1WA5m6DZ/OktfC4rBhJjiPjQ/C2D9H93m62UKsEB6fqw6z7afWK4glzJ
OVF0xfJsTXBqCsqXcL/9VWhVdHbwc4bzjjqLwybH3VkK3805rQdxjifvDJL3squkKhUzxDhvqxux
YCXZq6pd/HLpWxKlzPwFtZfleazpPOJ/L28rckt6nO8VJCOXJncTIoeCMgCAXuHqTuszYSZ835j/
ndM0X+4+taghccqD1JgV7Lhp2QC1mPe0lBpd0g1jI3+W+HiUwYstKCC/UBcRYBJpnXSGFj6PprnM
J11bjBcvjLi6Ep4A04xRofPq0vFjWX7MAvF3Okv0YKpYO/bqmIkWoTHcilT1AN+jSY+MdWlwLgxk
TmP6QwKTlyckOV2zlRNEf+jucS2Bkdeh2D/EQghSzCq8mj1DhPxhxknDNtdoAt/n9o+F8WhSiRfa
GLWeq6z0YybNc+5A7PpqHPbSv9s4YcM1jKsL1gEGjKV4w6OZQL3kFNerCQF+q2KOkAJJIzAKW/Em
fZZu/oWePBfO5qfPaPBgQ+hjyCBDqE+vmDsZaQ/1Pbj9GaxTthNM1+zPVWGnkYK6XZhkNV4oBgEW
TYdOcY7FHH7byBJnkMDdWcXnWVI38BzP+ISKcQeSql1hWcn05Txq/Noht7uTRSOmZsdplNExUaCv
TvQYeoI0YDzo08nwbxyuhFZB7GpKNHXIFJdfHBL9ioxWsdYXhmaZci3KFVtWf3kHKb5XnJJBThph
7MY6sKFsP7F/Iaw0o63a4nVj55NobGZIFxFljSWuSsh4Icz3EzpwiDB9tyGswAy9Y5LEKWvAhHPI
zM1DD07Nxoesge343+PO+D6I4vBrej9QqhVIqynnfjJQ2Qmlytz8HKKddQ0CTsrWHtnNF+WH2RSN
3ey58vsoZiKthlA3WFzx99hkHrC+mVZrfvBcyqioht3wwtX11zIPsOK4HY/oMyyFaapjMb3iWRyt
/pwEXwGGVpmSuXOMXLyfapUh/FyAgJD07zx4inUdyIn4Qw3fd2C/0niRiEmf/NufeEGgCzlGLAiM
VClSSJcH99hVXQxk4VuigwEDfGvOJLLcHMRlpy8Q7mJP4NNzRsbXxf14qPTuqDVMuBht1hDqQWoE
HHf9c2h8XMrC7zhRrL6YMmHFwf1ty9ABywURJmQJJojumeo5ji3Lzkm8wEU8q8GbxrMzoJXAomio
IvjEuHxB5y4oDIjPdfQhhjRZkgq+Pm6u7TQqUylTKBR30B2T209iq3uzLuZRjD+GiiMD+adqXnBq
0rTfi3opKxK0xDN2GBJMAN8jRc1mah5z3UOCe/wAo6kWLzpfGgZxDmZWPm7e5XnJgxnL6A1oUCUb
58PLjNUTrl4BOrR1AgRAZJmXIWivP5FgFNwunIsMZ6C2jqmsnCpffMoXzkNklAueWBEQXAcgrMDA
tZso9F2XHeMlruWUs7wLPHllsO28D79iBVPbg6ioQDoizEz5U9GoAA6s2Zp6kzGy+OQKVXhm7MRG
CsNPTGGbq12P0/udnAXZlGs2ZC1Jy9xfZ9I6LWNjiFIurvtiRW173raLh3VEpW0RwiDUb2jlHvaU
zAV5b5PiMPPh7F9y/d53fA7PCTIwnVDyj7OrolT2AJQI+fzZnQgH/8+pwqBNUExnGRuMkLYd/wNm
JhkUPM9P2lgj0Ql6+SYNsllzynbXbwJnwhN0CnZA5IOGWs7CvwlZwwW400TcsO3wc6LkoR660obb
vX+JOm1prj7/A4x4Ds9q6IturUNP9l7jx8opRppFDTsPc6/pUk9U1+HV/+0PqfB+Irivj0qvY5gs
eIU/nBsW8Hlefgi408TcyX+c8ffjhg2714Bk96q9X0OPiRTtQRDQnLX+WNjIXkuG2S52CoHY+nQt
gdQ2jSHKjGL/vvvAcoTzb8YDDe+qVpywkb4LWxEzoxiV6Oi2iKF81lmY5T2bOj4SXBRfPOsouUvX
lw9bN4oowXPqhwNvp+bt/Pm2RHjdvpsm+2kx6+RosdjLlf+7/XZVcrvFraFZ0EOLp1wJLNH6chMS
3hrAUhRxM/SeEmDlfIguM+33rL5H9aSUMmrmHxlxOuWVGoUH3DItCLc2tdXyipYNcx6U6Q7buTGY
elpN7S3wHKVwRNOHw2VMA84qsivowN6mJM9TrFea8EyAVDIJb6voyLcDvlSk4ExgcrPoPILvoXCy
A045fi9jEkSBSzfmWjY02AJi4E/L/DHZWT+S2rwMonptMWDVkA3XnlxgK3bqwkrOWFZpTQUNs2DN
79YHI+FUUEkduPvlleojDzM/IOmjWiQ9QV9xyS/YItLX4HnxkcCmvr8C9vrKEq3M1y2v6Rrltkpp
sgvWOR6RVFhGzxn9Ms56pvcMIIbZs/UbdgO1Du2kk0ZrLTcNa6DpE0yTXL1agx/9JVf2EXDRPbty
uzQ980QZKsnRVIgn+Pt+dFyW3f0LIXM2vG5T/iL8hakXfJgkika2S9Y9mKnr7pFnBfJT4KSg6N57
DOVcDA9VMheKjUi50uoRwIfJ0wXeLMtLidbRP1bhMTvHCXzrE3gTmzg/0DfU2ZG+e4Ql82IPt/qg
1T3RggelvMg/f1sYRTTPSKwevloczAKUvFoHKwDJnAXqOvf0k6U9U1NisTI3EugIcGQBQoNVOCMz
Xqnv4tzmleULvwMF+gDEdpKTsHbAO4MDtJxT+yOdB7mvqjWJgEBhn5YHCJdZDl3d6nuh7x/vzfkw
6+//HzUGL7NYgBb/RtKpG+elAF6e2We7KGaO1M95uVIx8cZPuFVQ8bCjHACpsrjuFz3ueVuS8bQ4
Pj3jaG8fWnidMCMWHLfb2mGCFi0iyRPn7nj8RssSYajh8zIZhwtS54jVutbSXLrpECFgGmXcqpZM
0uZxpAZm66JMG5Af3onvKGzF2tNks5QmbYfEBL+PslLInVYYSUdLb/Cuqmu+T59QlDJvOWQ6LjPJ
QwbLWhsGBs5X3k/VhSX9SV2g638tvHQzTZXBVmOYBgqAsdoXg/+vVJccSSpy+X9q2cwDQ9E5Ezqq
xCXe2SvhXxLqwAHmr0LFoOHyvQ21PWVbAfaC/z2ti4BkjEOMtSooo561UD47VZ6JMfHYG/C9vi7d
CNh0efaCcOcwtMvGRPsieoQD/iTDJsUsTeL68FRFoq6EXake/JDIuQxtipNp1B/mIwor5rvcY9VD
OuKSxVLJJGdpDRaxhPRmmkU7bRk+MggQo+ohBec7tHdeGjA75mh4XPqwaL/d3u1+IaOJ+Q3lmERm
lHNNnIHwcG8auVRP95VHKVHvuDNkT/LN1quZo4R4JuBB7ThooMgTgwdEruaQS7y2K0sTI7i802lv
tf69WDP/K3PGQOkMhtFkPJ3XYIL7V2PA8e8kBJw8AbvX9hSASJtP3Q5FlqeI6FTqoXh2bJa8CbGe
vnijrO5IszF9sAIjyuo1m9kNvM+T4xpvGbqSebLxtb1XyR0IZcyyWJ3TKwRQb8M57jGh0c310wup
W7ZhQWNYFtNY91Ym2iqCI10hMB17C4MdZBGdBOsXbOfN34hbLTU1qPZUWQbqA7YCbTT6oM5elPNm
Q5Z5khDlLAgMFi6M7lKlk9fVrjlTA3D27VgfoAVw7rF8GitgDKmR248LHbEbfA0fmiq2JNJy6GcM
g68xIRGJqYvJCclwsgjlI5tyLGQ+bRRUDzwBvWQf6dC437Z8LhJy+ZIg0rWaVqwhf3xI9Clv7fnq
tGxZn57Lbx3VW7c2H8qSZFY2QXlWJIPoW09c37Lr7ZiHpkpfbWf/OfpNG/PYoUNpkSbDfKMK6F7g
tPiLYlJWS7rIUHv5yuBMoqmiiCKG3iBdGC4xvtAy6z1GweWEgzDhj7bZQl3LJRZ81zVsZMWX0zuP
kg30Ce6yUmgQrEZLDtTURM/ykoIJCtlgb+gRm2al37YB4qPk+ZR1a+zapYILXixhjGvDpmUUU9iI
oyj74CZ0Qz6y675xQcBRsEpx49QVEc2WETUemIwkHsAiyyVlYe+4XrQ9soLkMTJA81qArehKA9qn
BYRvLbRMfQgkXDjwiWOqar8MZASwH88RP1VvWiSToZyvVg/qwDDntW1StCbTIIV8JXV9oXaMa/Pv
5jLDoM8VRjvijnazqJFUJXd1u8bKsXyJ0KR0mgPG4Y79sseAZgqL9ij5EWxxfZ/AsJgEi0us4CTT
V7O7MudF/rK0tDuRdjVQQQ+tanhuR/oqvm1ayXegwi3hda6B3vPty71+9OECTtdGOaIWebNYvwIy
Ej03U9WWq7ZxXk4sTpBUlQdnM4x+9hlGvE9taGdsvAU8GX+696SR+9ZLFUCNFWGCHPBI4S+Rd2es
eM4FpGECOHp5Ya35MzsUdyHJYbA3bj2LfKaYUh+PL1/U8RwaH9yDcDdqI2/GB7W1ZpisggZeHGB7
vaMVok8WNrHlRRJQvwsqOH4/oq8ouvt/I/EyGIFKVppqGK8JjPVGOEO7cP7tPlT4dnhOtfsSgN0f
5d1NeCCs0WSfxvQ7PDN+SNgYDO5TbfuGC4NA5BlATcRQ992+Qblu1KviXg6Xsbhma6hqkgzKIxxU
88k7egUgcRUQqpkWgbHb/6JKfTnqyBwOM2Let0+kwOxJUkkrvpQqniHYA2dI5qBoI/QSCuU4Ey4m
2+MQHTKVALYLNZ1eu6Ah9FJPc4cLfOPG7Nv4Z+FEezx5rOMwsFBCsauQk/DFdsFr2V2KBAZghkCh
wrunGM/dOKxEaoj4u2YKpWrznuASfp1yM1h3cOQJxaLCnxgdau3QORVpaZiu/HaszlcNm5I+hZ7n
NEYc/elnj7ggTPCRDCh0zJnwNHCvJprUcB22IY1z4HLTLq9N9hXHpUJFWt6r3mCmfIDgY2HdGepM
4fwYVGmDrBJVxRD2fDXVR69rnpV0K2zFZ3sgLNgxBscBRUxxN3Fpcv9dznrZNWr+GiBoYf+Yhwxu
hzranPlFzMBdg7+2axpaNYcyGIg30qMtMgWlMWpEMuLvcBoYSXWRMRA2uxxScyn4Nf4Ir13tE9SZ
V9CYSxNSeHvGV6UhLc7UDVcNDP+WyvY9fJWQL8wFQk4PWw3BrXdlGnwKqRZ90PMFXhHLuBbLEf7f
iEX3sFEaE1H5ZhJnPwzG03dw/SrU5tH5bhjLWh7njk4MEZRqZ9/3PoKrl2DLUh+DmMHWittH9js3
xCmaNZf1LLKGRVKwLcY3TViBZgpNHMAwbiE2u/j40soN6BlQd/Bb8GfHbNEsyRuPmiRvecOuGpKt
YIzv9H6akVBMFrb/FmUykKw10OL5ZzYE6gvVZJJrCeTa6t03lV0RuXhWvpaVkUdZcYaipPtYc95n
5C3CMKXhsAHKqptTIBCSLlCTyVQwCd7hDGlEd6ZFWVq5Y+tIW2xOPwaCVSLe4/MC5YWnvXLIXaUJ
vz2cmmtULnQGTb2NvzVMeAHSeAa/h/iaQp5I/FGBo1ARCLNtlgUQFJiZccxxeBOI+LJNj1uauXTB
oxscKvdQJVQIbDXrhczpKVOdutHz3My1m8K0AAxq0DTdLPRlrsYpC045vsGyu0n7faMzydrkBfnw
TlkM7Ly3WwKA9s6RrSUEzte8tBFJ5A6hnr+bKlRn1GZZrgo8/bpRtTMWoWzMN1dUM/etIawqFkDS
yAH5Du6ECiDtGmQo6g7E707ByzXUHgb/w7ag4zoe0z2IJ0ecqflfNyKc+18tX6onfD2O5hPUIMcm
kCqP+6P1QFx1ybhN3U0z50OhZUIGfl+cVYH7rugo715Qb9mY62LXDEmS1Hor8BKtQnpl6b5STYKL
i/LLVIA2CX8V/cxgD8oN47m/Y1+c7MRKNMxk6gH9PPFNs7vOD/CqZcmtUsDP3zfafhk8G6Q54fCN
OWxFcSI+wGYsy2/2rpZZdryOxuUXWAsSgt5BsebS3y+5rQT42f78uJkrCDd6QEWSNSE+WMgRzukq
UwxVmRJ8uooCMzdXeSlsZ6+4O/p9gnLm5Lx04+a898/fKtj7TTk28VPqEJps0a9qzpqXhGHOR7HD
MBljyl9pLkN2Ku6Xu2zG3Jaq8ThfJ6sQZ6/ROA+bSA4f7uxOEbNLKQp7gf6snzzFi8tgC1XL6Dyu
IMK8r3b/1ZX8WlqEf0pgNMY3gNlhtK3Z92sBzhkBS6XrLsMTVsgAjfSW7/SsNK+z8oiYvx+uiFWw
U/CgGNxDgLvZrKT5QddUulviXJfwRx/slwbAPEWcUpZ0y3qKrseSEbfZy36Yd82bNPqWWoq7/O8T
pAU9xdwbW0MFnwVZTxsqx+CJWtqKNArzy7z+T8j4lLPDFVJyKnU2vMqyqYR9dls1LNljPRXG8o6T
5gBlbD/tF7NeKAODFLHx4NSCqZgDiBV6W038MheR91787aliG/B54kNkHVbKpvuDyEnbdSlOlg0K
BRDphvWmOy4kfTfVFmaHQiuT9hsM/JMUqTNpIJMHTbU4X+JcsydmzkkCPVeSUFc/P3pmFZJOfn+O
rXgymC0as5bGaOQ4Gga91yCWUWGP6nsL5a4F/C/gcWptqvNFojI++nOUYkiIceirJw/7UoxjJlMo
pPwrwlMH2D1OWZF+HSy+mjKT2CZNWRVQA2dq9SLB37Wk67VU7G9VpdDFg765CVxVNJKiuBgfM2v/
uUCgsKB4zPALF1ydaRZSPCZSk8RlE+IcO6N5o53iSiZ76F58d0eWN2X9fzguB0PywwINoRHKQWBP
4bBH28/juae2Hgm40NuMvhqjkvXX6IvivOax9uS4/nWVh1xPAD2hbvij+1kwyVmA3V732fNRxAnd
e7Apkw9Jz/Nvptd2YdnZqPinhEJ2B9LKcoBuuQ8DRGuP6dGpM2SvjcBZIixAjxOFGgOwM7EgST2G
0KfyAXYmkT3ZpUutXzgSmRFKD90eW9Ah+TKKvUaF7AhuJvHxc4MUAr7cHfkBqxNIAMqWsdRTAFG1
A0wkAfUj75yM80IrAr1skXFtFoAsfKSQSvvIsuLlw7QVisHDfCq+kGrAwyXlYvPA5Yf+IxXk/c25
CQ2n394LaEBX05qz4bInRD+ETqFkRtTkpMJ8DCYf2JsvE07XZrDTMiHg9jlWRjEVgEHDWwQ2uVfK
e2TevQNyrgM/1Wevy+CpBnU8d6o55NgyGg9ZUtg3e1YUSJWXPCkZ/D5IGIf2aetaQphXlyozw+VR
1Y/PBRbRAjh/6a9SbJTAUF8pVU2KFblf9ClYB3SdsckU4Z1x3nnySr38p5q1mp/PxYPqidONLwfb
ZF+/OkAnW1kNTTJyBlIFftaXexZjkcY/jYRJtlOzSyb5NafQCmiBLzP3Pen/nPBn0oA9Mj8ozIyu
DVvFfoR4DFEbiIR1r97ViBpP88wluz0XWVGMi7Sc7rAHob1OYZ7fFUOvop0PJ2ftxT+hCUvo25ar
IJYylHANClf6w5eCzRhogGw0jounEz3Sf4d2ZaxVj4f1VAYhb2vhqrrKGlVAWJHeQiq40uxw5Tou
m+ZrxAwu4jz3DIxSG6Tn6ImUSOhcTHC/aawxGnSR6hWfQJPghqyIAqqIT5pFEoUo/VwJJ9sid28R
eLXLtvR6RJt7go6EXr2QYOMdqGzbyhy/Zyj6wfwjNcJ4HP02x1h4N1t+5omAAmEYlJbvNEMUDbPh
OyGbV5QPgajeBGjhN2kbMt6i4neGP3FsP7qW274LCq9amIMGisQG9GWdu+NyRZP96nqPW51x2u1Z
U+La7pGd3WHppaSOF+w51nIDX7Swj6yBHz1KmuJlYkQpQOVNqQnexDO35LzjTXmvrMsPluHzDuFB
uv6McYsKenvJTHzThYOgR2mNtYXzu0J+G55zrikSPHkeSN2ycvb50pDcgNN9sSIASW23BX3kDd9I
IerqTH0sEHx4Ht278qmlet5qBfWF/bf1gTl/21kLpBbZgHnMKz1V6MPmtMWtJ+DqLUMMZu1AXaCK
eSHx+Pbs/kHdH3f8FDT7yYg6QnjmeYq1m5iP0EvkcOQvP6rwNTHYuYsBNkpmUZ83/bDvhpvYOy2w
XOCDlErr2ebsJMgD/m8CPiSafDMELmUcdKRXdYg2pzMAquYh6n15EwYUOWWjXMsEJVQwx/DDkDiO
qJFhm9V1DpnUaOlcj4DvmSYCEMKDsCLcDQ7fW+mr+X4BNUZOBWbNnj1S1duAgRhmy7F1eywaH4dh
ECLVZUF7WgFNIPDIjTbrBieW+YlLH1k50J7J5q/Gr5R7Vhn3fuQoMdcK3Oqpncp2Qt9MZexl7rnv
GnoYyGXCswmG2HA7QoGwryPONlhHeaQFFhd/0aFPuPydDiQ/4DU4R8oajASFnxXnohYMh3UAX7Ws
6R3dRwG3M7zc6Lv7A0wBBi5v2LBbHILmQKMOUQsfM7Vr4dGsvKXAFYAj9c1TVHV9XISy89wyouUR
yTZPB7QlKTnQg+HvJh2rN2AvE773oiHAncAXq/UD2XhdOy6CSfdnn/MlFSOBEkFC4rorlN24I4QL
50ljUr9xrkaYNHw2mJMAAJZO00JQeldTPGpMuVnz/+8N9CJ8HN5zZ2x76WVJMbyv1z9Bse/h61qb
cGsOeeM1hUVxw2m63YkKPD7iwH79q8iV/Yp73DqhFonhj5iAnHEvBGUvYCziZ9D8E2qQFVC2AzFO
v+d/cq5JupQ4b5Hr4tJNQDUFumV5Wi5F2ha87uMZdeGomm/oQO+Z6UKcWfCSCraW3gwz9aakPX50
zXqMUEBTP33peesmUdhNnVr8+B8EhyuW+bxxsn0D284uyTtuy2+DF+fnCD9QWPdRIWZg0pZzMM6d
H/nmtCbHAUUlQg6YkLaG4KP0dp1LjJw0/z9zlZiohDuj+XiRQCm7rWlIjWlAUKG7hWpL2uipLNmS
SYvilB2HZ3JLnrcAX+NmD5q42pATQbiLNb5I6flUPWYi+B1FRNbZcPC4qUYsQW6r7PX6jgTdTctg
sMa4gP3iLLRmJGwwruf6atVz14aWvvDpsnz07OYPR9b2TdVydjfv+2PUuwUfx9b+ZkjYNrAsTq1J
acC2pd+9mRuSRe+QWRh9RhpkYjhAu/+64rSQ/TTR2t60Ege8WN19K5W8r/vk/Hc/63XH1szIK8ym
9staGN5G7gucuwyQ7a0jbQm/1p62mYxXqxjwK26ss4ZkX9qmiOe37ikQ0VPSLGgs+NMSHwxLvr3g
iOgQVOYI1fncrvi9Gypdrg4yWLrFYhcIF0dg5Al2qmMCE69F12UpV7OPfMkCNXw34F/hE/TgZ4Sr
nG121JtJILVQrGOnrdDI2mf+se3z4VwiXbpHiyYaQFLywMlPCa8PSrUMxC0kEidKbytQn3LCdvxX
71RdQ5VNMUFh9MYzsGsTqoiBAh2kozDPN179v5v8daKgK3f79J9C7sFUJPP7UknJKLSlQjH0W7Z9
cgNxoxLZNYkQ+dDOJv1szIIn7rFfGEG8/AF/iuV6D5R9GR7Q0pXzMpIs8Cy7U8TeN5RF4groqb3y
JE/G+iD4lRI33haCdCIwmF8aXf9YevemnMIcw3kmpVjSoL6It24gR60cCytGTr6n0wLAzN7Vr7tS
cq1EXUznWmKxJk4B74jzhIUKO748rAnpidGQz/9Iwuku+nJDI40rXkZjD+r0ZqoBJCTVidqpQA2s
toIXJVO+oThsJDBqhX1Ll2fFymjzVkMQkamDFoZ5BZxdwCik+DUPpEbJlEXuK0FN4syIA1QlJEkv
jB0c96VNSwotOIDlcPhMmGBurvtgK4VdAG66+mmleVdqe0Iv8gwp1SOgw9FrAzrmte55P69VGOVS
56LC5aeiBZbxyJbu+uSj7rrfNaNwOolGCY1JuDkCXcnGTIzl8oSRgZkY6WgxJthz12Q3zbm4BXTK
h4Lr3dN/VURdJN3ej6FPiXDDScszv3rczXEy0DIfJUeNHEIZrLPCnZnh3MQyGSKgcMf3ALMUjHjJ
PLf1FcNBtTMCTbQIS2i93uRGn7vcLNDzaGaWL0TtAkJDV9K1w/9m3yQnotjPeOQ4h0lG3c5OyVSp
e9tsJndXr6bIB3eyTwyDSZz3Z6Enou9KopjJOmdjzV0uATSzPFwseBd/pS4bn3wlvUXUSPe4fSbc
lMhwObKC4BpG5WgK41yb2nOnYb39D5jziOz5dRQehsjlcilfFytgzFUqD0K12Yp3pWLhEGV+Lfqo
hvvwaRrTC6TP3RucAXhBW5mWF3J/D5v8mx3Yp91JuFUomFrjAb7tVt5dGsmzj+ewNhNF4karK3yi
emncsGn9gT1xhjqsW4x/0acTPBZWqmxGgPUt931a+bKjRaLFNVDgJoczq2BwcldrhhdFNpVpMn61
Cyyc4c0RPICreGw8k1849EmxA4FSET54jmqKANYWH72OgXJutbJbgCn4tfEhO7fdv9265+A8r0qV
NW/4uyXkqScOmSIIEJuE7Hpluhi7FVIG66Vzd+2qk2QcfE9TMpCdDoDr8dFySnInN9GY/Y2gFCOX
ILlO76cRwcf8MVz7A0Gb7nY5Q058vqGD3MsHPZNK41lyPvl69UOxb9TDOt7O/fZxw9gL5ldCQdHs
yweb9dB+7wZO2eg4nKjqOiWZslXLm5OUKAn1dIhpl9eXWSK3FjjbPqBcXOyAB3SZ8rAWdMxM7dJO
JbZB3ex4EjXzIm3Q1GX2RkynXjIF0ojQrzDOaKdiUIt/n1zwhwEjhOGlIqrlqlTmKOH6DQnmUCoT
/d4ntnbIkWMbuPYXy4rqGmuyaOtwBFTzTmivwpDAfJcKm/y90vUcAcqFQ1h1e/RAxCEzf53p4m35
U3c3uXXvEDUT7X2kWGhKX1R+mAV6p6rudhGoNWKoidxvIsr9WhUFCMdfp02gVjSYI6uFKrDRfsCm
kJzCW1sb4G0TjpISiKRMs7y/X+k8jYF7tsPKuFQbgObeeVAxV/8jkWsH3ilJ+JRedzJHzI/r1GBy
YdPiBxiy9rS85GKR2LQxvKRo9h1sttq01xmzPvr5CjnoAKVoEnqX8W0bGwUn/JzI9PkjOX2+zkwi
hg3LcQCszvZsn3Zce5YkTOAoRlHGIpVRHGDOP5HcuSYdBp6r4909dX2G0GiSZjXip1/n4kQQhhF0
inU7ovVp6r5i9HWGPLAOKgDSkDhCM3ARrzbdmUsFsK9S/hS+L2kxouug+siDqTZWtVpUn3J9o/0L
/zzyl6z+7K9FTQ+4qzwEsUiUeA/50XJHV4eJZmxWJ40UmoKt975Lsda9ZuO/vFqDKAixXjqqDax2
lgl0H5wPTi+t7sIYHkirawfIsNQA+alBDDOa048A99QgkQJdOmeW+q/D2NI6Nof331+tZ0h4B+PH
NKpF3BithRjuIAfIjSdMhku4CNOHc9WzsyEhNwj//OKHIygvPx6tgoETS8n4WHXoc0QQKxnmiSjp
LZACHiodflsOlNsvVXlpmd9bneLd95kRhhBwztsSB82lE66i1xoSzFPLi0nluAGDFDfhMYino7im
MFrfMnMZ9CaaileO650tdB76sfSSpQQwiM4VepV00MHhgX8Oo8SBf3yEhesbG/YllL22cVX8SyAr
woGw47E7zN6tz5W2B7wQJup9fX6HOn0rF3zuP9tX0eOV2OyZwGR9QgAi2vgYH/EsFh+nc6GhQ1fG
7erGs2cVShmEdbEEBnH0yBH/snWVnz5LKernsnggzo0waKJPOC8Ms+HL9si1dGnA4jrOocaeJJQQ
tmaizzbXPrp2HMKj/pXmeOJHs1ZLCF3qT+heUg3PoX2RRxYl8G8w0xkU+iZAbRMesHYAU93tBGxn
3gfSALa/QjrZlU8YSYbQfD643e1JMJSD17PgEJpaSgw2zlth6BG/XOSXzYEmL/kXDM05zdjfP6Io
3555NxaLJ4Eq0FJuOubMYk/nyFH37byE/5d47FPLF+NSlmwkPwgfaa3DsX7tQ1gkBU+2L+N4+Gih
EwWOI3ZPHVwRWYJwhXUKg4CQ7h5iIXjr7wm7zzrBVDL+sHKPP+GV3q1ua9uZdYTizGr3M8FoNcSM
LDBnAYWyKSBsT49MJ2giZVzVHCXP5pCo4mnMrW7Y42V6Ka93jVeQ+Ep9PUQoth4vtscQL4o9zsci
Ah8UXPs3FYhLFM1wnVSy2gY48VTNtq1VBp6jwp0PW/LxzI8awJnVhXvmkmU4bc9Uraj3EMH7KeXC
wG69NHycR3p0tjrKYiueNO3Z5ZZZEv50Ex1vNxNIRetL5cg6y4HPj2dwKUmozowWjRfwjPJZ4JK2
c/qoy5HhN0lJ2IcuoT3UhxlHgZ2qpjBbfZUJssX06HKGV9cegQcbAQuQ6qIU0JoT0ORyXeEK8N7j
BuOr2/V2xcr61XkfsNFlTyjOqzTSicZVG7aDkzZFXBRTtXg1e1NHtneNxdmvyUmNyuJm521qlUI4
yamg/Jmx3g3oSfRyPtdDt8Xxj+R0mSQA6siFKFPkI82WdAjff0GB/k6mNrX53I+1uLgOfzVCjkSj
HRUHnqxJA634GQX7PPQmntl0JaQrFACTXn3QsGrcrFwK8HrFnnZ+IJJTqVsuPEkvKIbZ+d1eznt5
zFEzIO4A+I/4FE9TC5/pG2BG4cfwo/6TjsIDSkZPkaXsqgHf8K5yqyB2Pgtsua2VSuAHhkZsd8iW
jollpN6et39VMUTrmi2T3WbM7v9Y5W/zR+dHHNubHHlMb2/t7zuQOPKsTA1rZDOeTC0XUgwAPBhF
GjHG+vl5S6A1hgXP5ryjwOAcsB/twwdB74/oUpg5y5It+dWM0lzL0EvpapC6+3YgHjnQh+GI+t20
XfF04Ew4RTwsh1oyHQ1Rv85p0kMSlTtGq/UPnYEr/vtA0leeo6JG6iIoohBHjEHfRwQHSqOofl+3
JoNznkvdgveYlN5wSuxxjRJ3FN7wPNLb3+Y3+yKkM+1evLIKpZrHUBvA9Jz0Jj3OK2ifou6N9WCR
J7525lAZWhTJF1F3M20JhD41QQU3d1XZTfQR1yJaKdCKCP7C1W+dwNX3qvJ7rVZUDz7tW9lUr0g+
lTfUrfKacKuGBGMM2BIeVYqGu7JggSTxLmk40wWJzC8SmCVjkCXTloQvhfwm9kBuIncbIFf9OLV4
35+OoppRQ2q4fvBHBkmuSWFcGziKjr9OF3TLMIw4mhZQvX6AvHwj+L67ypBNVEdxK1AJkdD4QwOT
cXUHQqrzBp4lMxaCDfnHPkjndNWzOc0Y73SQjTTYrleLCRQEhvnCtKurd1uOdaQkXIhlfLOrxa9P
4WqplfRr6if2KW+ImTNbOm/40zvmBjGwcO7oG0MRl+4twMbO+Eewo1/5vCzkytueGvQNzNzU2FNP
sD2EJRlk8/YxuYiPy12xgiEH+dFoaqx3uoa+S9NbqotsafyoXc5NMPRFmvuCubOdJBIbABCZt/Xj
tyHyYVbr0SJ4b25g5D1UTfZV9/fmuo00WyxkPzYeY3Pk/dOcR+0eNVhWyQVw4ruO1DkroAOzhcW4
nbPVIO/9njebJ6yuvr/VFGJgXFxc0zr4paSDP4LRiWQILAp/BAgbNQn0zYsQDpj8LfPucGgGg4SE
WQ6DevNVfOTAaj7XD6Oy8B7R3cPilGm0VMnGV/sjbSixB2M7wMc5ksNJ9bKbrq3fQw3Da9ZtgJvN
Ls2ER5mUKbafVDF/S5xkzMbJc0wNozk0sv6HdGVefQ0eKYxGqUcmsRFwGkZSfO2FieewyRZPPYPS
KBOc/hKXaZY1u5ZShnYj+Wv8aHaIe2RGdGMdXUvZzwymAwf6Z4Sl0Tzk1sKn7XyxX/V9jugWQMTi
PHLPp/rfOhENBqO92UT6VfIf2kkYRdl01xk62DyDVaZVP1Z+z34mdPkZm8NqWcW5mU8vPym2F07f
hPVe782aPWkHDCPtzDpnJRIQTAd4wF5cAaJmuJjo2yi2ZMCeVh4EL3fqiqvT1Uri+Wq7wtxHsxjn
f+fxfgjXnB0mM+EM7v6wRkpOH6K+sEkjlgdX/9UZzpiMixtqG6K+BdS+zZN+E5b6dn1FLrZwMgfg
4gJpXdP2j13dumS9buP1oAx2i1+QBoBg+S15dMioGuGFLdtvzCTEZvdooH05gVvsyOq210OWfmW5
fiohenln6UmcRqE3tpfGubh1He6/YR18Tm8ozc2kndPDENe3kQe4ex9YDgr/caYZmyDXkH2FCOYP
SZP9i5I1vsuK9mcI5S4Nya5DT0BM/BGaQJ8zqTVvMlIeFk9YAXO2lUP7mNyBVz7V4e4UNT5U8zds
XsB5K8f8YnjJi+yLfRMA2n1etgBiqnhAZrqx4XQJc3f563S2ptJUGsmkbpr0epTo4dMnMzTE2hLB
IU9myTfSurc11LSakbObvm2qi7S18WjqkqCIHAYoGe1Y56fCwA+JVfa/VJ9dwzKImAaDWStmaJlC
MMMA+5LMbT+5dGF22RVzkBXuc3v2qF6VIc4YZg8Ilxx6M1J/8y+5q67I6zgxJR/nJa28S6eTHsV3
0JlFMRMyY5GE3gQpOrSQHSRXZJv223944G4Z8OYSwqcnuPxx25tW8h6j+i/CUEKLkfb266XMsM1Q
+6jMFBFUyewEpnRoil2SZFqTomnTEPiuj65apgyWdyzF7xr5F63/jBWAcLjEzI3JjjjOoXbWtv7d
97nwazBSa60r6soqU1mIpHiltwby3vcIYPXOasbSE/d0E56flQbD4jtgZddHw/O9yODR+gvDgjAq
NPAwJd7FH0ebcO8Rv+LnlfVkr0sG0fC+sgyrmb7KyF6x2OPY6WF5i4iNQZzIASf6GjKEILTc6YvX
Y+6OtSjLlu4gCxenv4Ynn88zDHgZsqVRoTYZzGkQiWAzwxV87iHcqhDrx1VeTexz7YZFkzrDthGc
+Z1VcGlR5InyF0Gv8BBrGImj2535HlnePmPmx9eOlXG9lYxgkGdC/PxqpcW4AnOjAsoPnnCg8DbS
vxTiEDnkfaXNldDwETHTVjeKLdi1Y+cH8IY4NCUJJoTJpka5D41Gmoz0pFbG9bHj4FYiZBafnfUe
TAh0a6lERlehmzKtZOQP18qFETI8Lb+9jpyvcYSyfTlFTrU6f7+RIx3c/HzaCP1+2s8iOn8jSTRH
lY3DjEmOsCDSV3yxukYVX2wzJDpVVBc8c18l85QR6OhxURHP+HvREpAjyamwAuAaIsytGs4yTRhd
521FLpKhGcKrDSgTEfBTT6de8uOArxe7BuJuwaT+tNbTpczjTGgfcXmoVncBS58fC9L9S/FxFSX+
cDrz39jMUn1ywaUsLtpyJACALGkEuArHz20mY3Q9R501NXpHGstCYo4YIKK/0FLh9xQoORO0R9a1
Eo/9cyuwlEcjmnAyQABRP8sJtSfINW+v7N8fX/aqo05n5WwBpueTtU+p+aujgl+vytHxxKNwrcLN
LA/TUPeiAM4V5wBQQUDlgllLYBV/VM0sXoB6Y5rC/4A3O5yojrAYZLFon0bAxNm0afXAPbw0GulM
YIVpvFcCnKAbK2/bcbRg3UVvCqvMqhkWtjFUguCXbJzKrgqU3+Xi6oWsvAplrDiXMu0z4NdFBoH7
y9cVGVDRadZ1FwFgXkwdPNtxckvhnj9RaF0CwmEbXJAirJOIKmu23Gd3zYqSdiKgSxXUksl+Fiax
M5yk1pjb5/z49RSx9iQxPnSX4FRyYyfPND5YJReVBi5NkJoji7hyPpN5XN0wRi6PirxfjB8mg9hs
NvCmjOOA52RXwFhAAUAVTs5qsONzIR7CtCYxQiYdZTej7aWmw+taKhGGuNaMuoaXAbFR/wsfCP3S
RbP27HyhhrGZ/75py36f4e/rpQ2T325kW7ucmhRO3qyEuifYCmVlOpMyHmZ/x3BPbqYJxHuJ42Jy
Ec+2zxdg0/Alra1GbAso5H3X4t0Wsh+hnCPOF2R0gTDQWGdTfm6xTL/u3Ts9yFWBLDyMJsL1NDn8
Zbk+xtLeRMRMONB6fT28IHE7i4IU3DdgFbHrgSsSOOPgyy/Y5hU1I/Pi4QxAKKdL4N7x1H3Qt3Ru
EqDvfslyVOBLY9E38EZPwuhTNUGCyPYKhT6R7fCEJBao/NJa8/PhXqf5ZQevSuJ2wpOt8g448Qnx
HBRQdjBKlpmukC1q8pnNzkG1V7F+k0DWbEuugy+Gwy4+91lys6c1GXp9KEIQb5GPBDJoPaYwm+Iv
+zJewPPEexuQT5aMyj/A/dl7R3Z77hZMJW6kipTH4gubm5cjIWlM72ylib0VmsbhkVfrA5n4Me/9
08DcNm7GHo/ecqcKBybfLzR4NGuIC59ZjftEiYd5un31zrtqfVCChi6E7PfsRfnydezV1Pc8F7tO
WE0X+y/NYGPsiUqTNiJzmw4CrWBEQh4kmfn7oSBUJBm7XhQu1NuSF3ESnBqZ2WXFKx6SzEyR2Y4X
LDg1Np+vUhM+IjpH5nJ3/APHGRR0sA1DY0jHGT1l6RbK9pHjSnzA/W03xU8wphV2+gN64CosXWaf
WmvIdQrCiV4KnKwP28WCO6HidoW55LQwTAE65sKfg6DoE7dTB46XPkjy1dlXatDUmWlQUNYDJMQa
O9DUIynDVi4ojzKmGkOaaB66Kh3zsdeDLHdjMP0qM5VSiCSEj40vjcDQg0W1CkqW3fgfm+tPcjkG
EMUgruZaSKU3KJCLGiVpwQemJ5LiY47HlSDcg+AfQ2gvC6MtZI8SqrOmK7msAyBQ7d7RgDoPkuPU
V+psi7TGl8JlSJ1T3eH/vN1DjYp8Jn6Gln69ppPOFT5LKysyo71zivYOCIWEfcdaDlYHQQSBb0HM
/2sW4i0yuE1LANEHWOfd4PBGOIPMvf89FyX57vKJHn1Zo6PGiHdJI+wJWibH7dmz0cTm2Ipx/dcs
2ONKzwYL8HJkaIZfxGc96iats5dkLqvloWIlaUMx0RLuWw/Oi0ADFZCcdlVgKZdOSRQu7NPSXJUK
6n80mMgIV/pegUySNxHhFmUGDPC8D+kfVtMWVTBeoqvuWyFmNXC1nm4PsEMZ5VoZAMrhmcP/JUAr
AKgmv53HGW7X94caoJkmoFhuBrEDwtkMsRCIKZCe+CzSOUrZ8kvCLPE8igcEdoyizUO+1k33vmaM
zRg5a45lGJ4wuQGcEtw6zZtpeUvSFSSdyXapneqgpLEh+N6GtbR95/Wnr5iiaEMCHS0+5EgkC8A+
Na1DSBMgKzd9xm2NBJO2p0TlxFQCXhYTgOUh1Xw9VkT0o0Kdq8H1NumoWmLn/upsUAQ1a4mwkJR7
drP1+7WvFqImyWdePpfCqAC0wGYli3LvhqwPKxzJLy5yrAUE+y2Mhle2LC9qjCQ71UFsRMxKVs7O
9ul44Y+D3o4kg9gvrmPGG7cYivVOPwYrCeGVYV6Hd2tFayeKpRJdWokqEILL3serUOh8D4CR2r8+
AMAWKt4vlCpOdrrgglaO9IuzI/idGIyAoD1VbwWzvTEJ8Tu6q2++Qmjq31d4BnXYALtMse4VfFBZ
+gQOAWPOz6c6p1BVmRVu4dCXGgfSkAoUaHGR2yWQXUJWhBRtku3cEA7/ZTBDtLp7xyu/2WlAOdr5
l82nYfCTKOTR1Lh3KQHQMLiJoppjUo27aGC9hn3kNhDHFIE54nn0G20WDiu+9f2i3CFnXOHMT1UN
63KDLV/JIE1a22YXmQ/+T66plc/AJmVAYfnn9xAQUZmDavUMHOxNL3xDWP91PZY7D6swxiMUpZJG
5QoAiWfAeaWEFHe1emVNdNspqsaWOoorRybmKKWdTCuoLZ53OryYU9Bzc4jJej3fcZ0jYwDozSPL
VY4Kog+iVjiV7AsXYoCeRmGja+EUqSF8RDZ51Hy8bes7+wpu5tS7JoVINdao3j2mBtdlWBV21hnF
Gt5wTSkurJxUFn1G/5eFgE16qB7Kw276NfL9dOXsq4w1w/bTqNTj8ex8i1T7JihcREu8iWp865Gw
o1C62Jb/VFHRbYi+QKDsLLaeQCAgJyB2v3ntKM8eKbpfn97MS6ZzFown15alrLkCXD/iUZ4gdOZj
Xh9EiF8/m3/pSK8EyOTdfRH1D14nGctF4acJ+nu6kRrRU9hIDF5SZsfcZhrBJjsBoC0RnQjuuDso
5Yuff7La3JRp3mXGo6ZyC3pNsSku5Ul/BmLVkUIgxA+Aj4dXI9S7+lzT79jg6fdd3nOQWyOUQI4k
OJqCac6zuZvFKVuiMo8AvAigh31IdV7phaamgBgEB8oJTReW/Bs1Ky59RMsg8dSGl+dRefCeLnSi
BlWtaSZulquVkG/476eKUyO7KKVwlOn05Cy7DKdk4upPmpCAa/VRK3OxcwGyK/yoXe0HjTujLlcx
r39+mPbPRE7JhdARk2cfxig+T11gcusxgA0MyXH4Tdlec+zK4bKYeXDHgYT1xcVF9dZVDM3OtjZF
tMq998swwh1U+gW/Fc97aRG32MeLXt8Huk1ZZirHJrxdsF+iFKgDwQPKgPvhq0RBVAfAQWJJQVph
4PKd2sBDBZBP7FWICfdW3RsLeH95LhMGd7Xr5oIsLC7pOuT/lCJW7XlmVXC5xceNdSogKoXWwKtj
Jl5kS6FqkHBZPX9PA3Z9w8S03WisLZHp3e8m+Ia0DKULkxZB793R9u40eyobf8JfdMvEujGxGf3C
q+JwZfNWpRQgXg5kUhC4X3REMC+RKsR7dCVO9DpSj0g/Qicembu5s2O+n7foIOY/BVHMqQ3Ou95a
FTmKIt3aTKx2VG/OGV7eEE3AUnlKVBBTl9Fpd+Gn5YPtZW1OmyWkj/BYO0H1DTYIqb6baAxY2WQM
patWiwuGNhK3ohHDRbdZGoC4HmiqcYMw2SOEZnnT0eipCmID0fIjIYaJQvf3ZGDUX1ROX95UcaIw
475/88Klmnr7ZACdeQ9OV0C9MRT5N9gi0cxfxu+bBpukUFOjjgkknbPBCqnOhA8NLMFTTzLofCWo
vF14GIDK4PPi5WIxXT0KD+dm/wx3XHN4Fkzo5gHAbicyo7YUy8zy2Rl547/KFu5MLD5EiDMm74m5
8dXL3O2VgvU97Mx5H+X587jlrLJQjV0n+MHnhD68bKrCql48xrCakq/4ZLZpZ8rkYQKwYWDPigvJ
E1xM3B81NI0WgR4Ig02mY/nkDcgN1G8G2qFHPS1phn2WSNryQOURmy7LQYJK5yyP3lTRCdcpb9zo
7Phs09WBa9GtJML4Hn9E8GschEVgrWFm4yatrmCavjhdF7u/bbXFN0FJdChuv9tH3qRmTvINH0lh
P6FXKrZjtHsgt7WYZPEyYbmsIu8G+ohd1ateSp5DcTGlHOQnj8f/vIZdKKvK1sz+u0CYN6PfsThI
Cuf/ltuxIeZ93cOCixXegcfaUUa48+wKepuSQAnP589cKwPEdO0wFkQGBBAW8zgntETx22nImM1T
w68BgbbxQkQtnr49r/PbKEF5IpsYwkgiG1cueK0hxTdEC+doGk7BFs8Jg5Bnl9AW+0pqkvEKPTZh
GREKaQo+63w68yRzu611avIE7p7ncpAeue2JKD1FggDMPIR7bppOhfvtMmLjncYBUtBY5Ts4up8u
e0DWlBOmWlB4bCjoIRnyRZvnaqzd30ohvNKUdHgNC8G2r9UTonUITYlm3V185ag6O2J1l72wTBWk
dgAPPMw8L8/6L/7dvQxb89oeZBmK9BVlF4gSyJRHUJfOdP2jGfJ7+cugQcc5dFvdpFTLvIqWlf3v
7wulY95jBgmI/p1qPM0enJeoPLgwJ+PtARPWKxszUSfLRjaSprXgjZGELiFFHaswsQDDAeoCcCYJ
W81zGjz4lZb9I7/keOUzHchwRVkdnOiZR76tnbUZEdfom0U4uF+goxIE3L6N1Vx+WNxJx8Ku2g7M
8zA4OvCDU++98seDz9FfZqZ+UCoYmBaNkiPjI1c1DHqzmWzaQI86Sy4kc0iTajUJdkyBOeV/zxHq
NOWol+8T1JU1Un8NV+vkbUVdPyk5XuysiiW4yH9sycwONqRLw6YUn4AuRs79Myq8qUzkWTBNkSt7
1ofXqhomXrZBp++uX+y+DQcfc0Ncc3aOIfk8jvqkP+ysT135j9sjN2K50pbNDV+mgd0yiASv1Y2X
mjsObqfXMqMZpBvk3dpkV3PETefMvpKJdsid9np9U9sjGdOBzsA6tbyYs/L87+pJaUFsaZciARoS
atfyiqC9YufhlQ4PaPiUOALKoeae0k0HigItoNEUkAqIHGUhx4Em/S5L8mDMZuX8/41prqnCHpSZ
Tt6ZGs9QwjdmBgrJ85cZP/ERLTMcYrtn5Oh1VmCKep5MCL47Jy5SAplBBLMhn0LvPQ1fDlCilhzy
1Lp3G7d4dtBB0NT4yv8a3NoTrOaONX9yLSJkwA8MqQsSVs4lNvLQPAu4Qbyq9oTpvwMgS92OSYVV
ebIQ1WgLgiW6NI1FLrSBhRLZVLy6Xm7Js10+kSDw9LQXclCylEvhqdH7HgtulthF+clr2+pe+yb4
DE5sRTsCMF/+DVWdRVw4Vs1DnNT/ASVRSJsbwqKyzEWcRo5lGxpz0sf4l+gendo99D28CqCN0Bav
/nYU11hvUPrY2xe3knvfJhvJH9DwnanEzEVzjf8NqW7GS7X5stP5ZY1TsNUiAGkFuJCNwjFxH6PG
VegeD1wn+M5F0s6Sy8CXilYdxG0HqHe6QJEm0iW8FakJ9PbZ7FzPlLHgI19aP8JnABCEl0GdPmSb
QXGkPlw8Num5l9aUA6yPZ//iLTtQ9ceRsX+7CNSdIS+WWHKfjAUbU4tNZYGPXlEtEUfsXJwKxXr2
+Trhg7ROo02/xOAxGvLkRvsZ144Vb03kZcEjwZ3WXbkaoUA4SaTjC18soNQCUfL5L0KYDqorlUxI
J2xOE2By0YEhNs2vgMw1wbSFxdPUaPGJ9+T1wQR/sirTClvkVxvAM8kPBJd8J5tc8IWRUxjhWyDB
U7ZoYiJkSenrLIsnWURmOlMywsqJjiImiZyp0s6OgGUsSh5FymvNA5UQaxR2fhIneQObDvTjdZWO
lqiTCnh/aq0/Iva+3eB8HZ/W/tUt/8WaG2EZsYkI8XPfPy5iCUlR0sbJcXooiWTNgk4rUSNs3MH7
6VoT3HM67TkgaJM2V1QE8mF8jvtQb3p987n9ijNt+hotqy3VY/3t1Di6TkDaNSVlX/gqzkcIq/N+
fDfAe8XbLFTBHNAsQe/RHFGWwQldGtQPQFdgozLt56zQqfQZ35+wTRRy2ZvkpDgvH0CMjGENFylX
tozWuwNNuCRtdN55wzlB/m5TTPAGuhXloESk6ta07Rt3L4jqy/VDRepQ02zDgFP3SdIK625QlvHA
2Q0/rV+rcAfvmMTE4AqLgC+Q47PlYsUn4JHBn2koJ2EHgrgGrExtgN0HYvrgrc6vj4Fx3ugEi2OB
5W0EQSXzQBMqlXBznlUIv6cAoGN+n5B1LYHWl/16gNxHX8ZZjwtfVjMAUKejYBpxshaccs2LGnP1
4PKLg9NgjirOG9TuCx6vW2dz4P0CaVXYK7Zy/uVBTSRq8sV8KzPcfWeu+cNmtccf/izGy8fcI0BY
j2kBviAB/0Cs+ZW7y0UQy6Z+OSh2h+nhguc1wr47ZNH//FtI1bC6Xb53obDMbRuxmzVvVElHuxpS
oN4lyn10BW8TKPqTF5rSZsBDv4E6/6FMWK/lIeqGCLtSNXyBMOLwo1Pkozx/8WO/UrnpPpbZ7aD/
zr+j17MZ2TgBPHODZqi8XQdtXgIi71sftHy1sEI7UcWOrl75OfQ8oQBE4H1q4mxGGZusv9cc3uXx
KMvT48WCoAtGQSJHektiiIPLNBK55pYqIuwMYrqqsupniKddEm2Phecei+2rSyYzheM7VnfgRdLn
BK+nGvkZXIv6h1vZ8Lfk20VF/jjCSfV9M96Zbj8rGyYTSR6cHlnOZYmD6XRw2/Ge9s0pAJLcnBmD
5KmaJ5EegxRaTv3ND0GkqjY0viPvylfumnh4wyadbvJ9Y6mGig7jB1AoT8wnVQxtd+y3cD9q8tzO
C+2zSVWGeiNWH72wCToM4BYJhe33UVkOd3cVjQf0adQEV/CwBMpVss8Fztq4NLDG7WO34iQBUqLL
1vi+6HmK8J2ffqiA5u7wAiGI2AHWo8zFE0dqXyeHkVw+NnxShBnsENvaNXMNtvKmuntWYGrv/LoZ
Qz6MBtFFu6lfxTwYgbCxrQUW7ZdWsYlqtsqEsWsfgniW+UBKXxDbp+EoTmlvCNz/7fAWjyBdOoJT
Jww/9P9wZddS69V3tWh2ruKzQISmjx1zqkWrT0oVFx9Ps0q7RWR05D5DMlrOWzyXIop/nFdb0y4d
SUrjmCyzgyy1uFJumA3Y1yyhr1U7u0Y+4JbXpb5mC8jONjG/s+y1OXiROvCkQj6zDXhG8nU5t+Z1
UOfTbnzuaBVVpasdm4QprosZ575w8yPOf0MtTLj5QYUctw11apZoMdgA3hVmoYCr/Fvjn+ENywm/
0/7zJXt4nW9+PCzOF4eDAlx5eW87AdruoO8Lhk8HJLovcMcOVn3IXxXuN5Su7urvH+9RBFeGRHVp
p6LVH5LwZ4WmNVRcbIcFIc3Z+04MqHA3YAbOxBiiRVOtPkZ6xFpPyH2fqrh0i/UcfjshLe6cNGF8
iKozxfHN93UyNNo/S9XulTpwBfSw7pkoxtpZByRI8HTMfq4wtiRpi+Poqb3iionfu8IUjwIhOEGz
YCT9jKedL8h3m9uqfz1BexI7Bmtck1avaB5itoKJIDOg6wH8n6MqrTRRsZ/tQWkjt+NuViHlHuBz
5ka9stNfBYsOwxgP3dpbn1i4DmRe8jfWUysqgI5bt0ug3soeTjI1KbEnlyGn3h8dYK2MgwU21HWr
LT1bmpC/PjkU5pxTIt0paFbAplyeAjEI6RXyn5Pj0wRNpD+KqGk9GE2dHdXBYN5++FWs0Hj21t0o
1rqsSzcH6jsu1lhSe97o4N6MHhdGezXbjMSNg7jK5m2ykiU02PAGoRno2zmdqCST2K5a2rgalBeV
fWulweegxXKlABOHBB5O3XjSz3l+WIRqZyAZpEaNqAdCZKt5h/c3C/FZsM/DuKb+Kph8XLMHcMJl
TWxLfS6lPmLZ08NqNGMRCpqAWCiIe65heAW+5rQVChKT70pU20V4XxB3kQ7606d8xGkridRFqt6k
2P0UYCsgIol44OMlr/DZjz5ZdNLhcYvYdAS92Xdms6faX+5JzPtHV+fsIItEZF1GhOgz+Fp6NN6A
P0dRwW0q2Hquf4yroRQZhsRhNkrQp3Hm+WvlyDKi3FlyEMUSsHcPtU7CIFxobQVV/XMNDUG4kDvl
szr5sZgLM3hRTnh215hKUGMbr/xdlZyfItjNFScDXWoMi74H7OCVCV/DKGDnh/00GkC261sejGAV
8vmn07r1DRFtrIkXZgyZrggX0rURFyDhlE6jivUPNmT5HSoYeenbTs+3VpUYq0SzeQ4rFYWqqN7r
ehtvVNFHRBxK2ZDYkFsGXxvNcPRUnKPejqTS4F2m5pZOLFXaktyQNrR4T/Lvbp/59pr14vRt4E9I
j2aOYrI5RI5FvQrvewzWZyEFsQr5WQVv/RFrplAnnu3jW0AlDd7n4FIoIqQEBJMW65zxKWsxhjTU
c2N4ZhP3athEGv+BGduMblNayh4MN5VaaYydxxsZGttpj9c9zMO/qdYGEOO0czyKnOV8whWYoHWZ
uivGtAb3H6tCXtX5RxRDuq/2vK2eiei5zsRTEXZK4osLDoKTyvzDrrfQGCVwN4/eH2k7iHI5RBay
NahWArB1z2AsYCUehU+y1ClxwVi762ROQvUfG3CPwbix0NzU720RqRMrR/h2cXvtCVe8RpsxiB1P
jv0AX68Pw5T/4ZhdKKkcncw+xBR/Cf3QQU64h9Z17j05ImbBIfEBDYdJQx5rrPHz2n1wvqaM0bHw
tQc/PtlxRhWummB5nQeYf3O/U3dG4KzsMI6LQZt2cM+L5fJ1kKvXMxf5rPL6aeHaG9sBU7BBemj1
9uk4poRa2kWv9y8i7sWD/5yuWc2eE0ouuyzCHCVmeRvP0IdezHp/RvyH0Pbzxx6oiTaW8MWyQn9I
+megYvOYDY+FByTU/OuaCo6zz7QHykCV6EO1h+NgiiEYUgnOzd0nvf4kDEag95+126U22p+zag5k
c4JGl198sXmpNgceiM6Mvffj5oK3bGX9E1UuYqVE7RHSGnv0kwog75Pp8lpuJIAbAw2M61kvgPCM
6m9fqDDKrNyM/o8+3bEs9AbiIfBTDvqktBHliS7A25bhTj21loWoOpsCioOZEfKYkG/ipTHa67qT
T0gALOvj3qhCLNkcNkUV5l/bgofNHWSHK7GBZuz4I7QD3FsMZpi8Lp+qK6rD7iNvOpXvOHnuUwCp
iQBiIga7OhJ8Bbf5s5iOz21MsxV/On7bLnT+DDkY6SRgiv7ciehQGhqPuwnuVTBaf5Y7E3BbRNt1
y0uXqaLKVod5tbz86d8uMAqxoADaUliuF9hDRqZy1SsYm8SnkjkOfqYNgdYuhH083dNvrDqUuRPU
1DDtMwuDidYxAYiRpo05VkIElZl0Gt1D51GHm3oBMRXEaPgYbV4fkGkGxHScOYpGuS2RctdWjSy1
UL7qJwy1/V1yPO85HjfvMZfT79WkkeT0cy5EPGiXYrHLoHkxeH0/v+yjpOWDlrtec/UDZVGRTqLA
2gMfiY3l8pfK6KWipxpb5sstI4nl72yK1fTCje5Zgf9sbda0zgtGYD6BtmU0iEtUm5I83SxxBUQP
6VRk8DmqsQ8U15wl0AR5HrGXwZ2fVMXz1m9EyQ42Mmodfqs8htUGnv+yIicKLI5NfIx5uhFlzqGN
vu1OW2b1IHetkfh7TtMlfodiW1P0LzZx0AoCzb9MoQAi3Pcuu1G492oeFpKeDNklkskkZEHfn6Oc
3Um7b37U1Y7XPxOoriEh5pXHydAumv/n1SBiauK04U3xq5Ia355hn0UsmcKZ3RXfV1JSXD3+jvED
/f++DB2xpV//YQxGcHldsrALFaWQsJCiEGzlqLEeSwB1A41awB3I2dNsyzPKZrt5ijSf+1i2XbE9
gUgOjcD3H7j2z8g/W6UnnzWRFt9voE1sWkMPQ0jkWxsXZNMyAjhcJPSDAnluIQSZc5Tih0KtNxZg
j53XMnDKy16rydQLErbHCOWoKVt8CciRlAn73oaOUUSJMpYEjaIeaf7PiV4E+/+d1KYN6bJcoiJD
dy4m6RCngNA2nsQM38sTQ1z6qiQ7zGGOZ2wXBHJ4c/MwwUp4BeNUs7Q8JvSPnXUIIIx+RzQtCzWK
qmoYPvoklS/1bVMqaxlK58+VAupgmfBIBfSayK2taWeSBladYbnt8Ye87dd7LIwKtgrojNjX/NT9
TkE4Mdds/ixMt2ZHEempxTNX08HiYnnyaEKR/qJM7GSyHt3ZYEoXHmWq2keujQepSZgkVgm2gsVB
KTtjW30BmrJE73A8r+iL5k77NQmHMZY9ohBQruGMDkqcOwzlQ9BKEZi+5wE2JXwE3dYdLyCd7sHI
dEoKWoFT7Cuw5YmeFi9YfPKqdvcjTyS7rRSFalqxolxG7cufkFQl1gSQfp8JfoImdHLPQLGojOn/
pmydMVvRUGXnSEXrpq5axbFUMCaMd/fn/AqF3hDt+KJkLdDqsl8UUbO6yHBUq5mc+17w2OeyyHIx
C9VjJZypvlW2tcBx3RuYfrMKemeFFxSf5Sqtiel4eqF9s8u2JFYpAlogvfqXVDymcyCofpfNyxW2
OR8PsPIRc359nKjgxKw3CRRuu9/RGUrKTI41AEqR33Dm+D02OcH+Y1Ng7fodYStSUg3CLLHO/HVu
b4nUIELkYnkfq1P3z/95s1s5FtrBOwc23v+17sneuf+CrhO5zlgIdyFs79eJYaE6ZGZ56JrUTn6a
Q5GsyZhDm7YVpW9jPT8HSZsg2CrPL/9x33nNe3MYzwg+LdDO81cAdq6xyjJ2wnjfXb0XqwqJhvtb
m2lo8Eq2Wm5GZr8jwm6nqZLSjFz1u38izpUS5LlO6yjoAohxeC1aDkgdcg/uDNCZFKoTHU7hwAJt
sa3wKL356agU2hW+bmSVvVr2qmMKeFWVNKchSa0Wi7OlYtlVphdxnHGrvsOkQyMtMB55zlt9x8GW
dX2xkP1RHC6vCd3DpVBDo/kOlsxALFdPqp+/TzbEZXywmZHaPl38Cb/mGj1rD/lo1HE+xif/zPkV
vEIYPWMq7R1Jo44Cr+pJU2X4sQMW/NtbjJ3e0VOHlFsD6hgLLI6j9Apgi4CXrnvd2oaDzl+QtdNj
f7A2h68/vmyfmN/KE6szevNnmDupC+xMvWl/5LZQWMHvUhPiGameWKynRJebeYdCugdhfpJb+rN/
IrPRn+sA1HgMlQoATju8XQS2/WE8LjSgPHOGmEigVDb1Q2g0AUrLVXqWn7CWv2brWa0AmXPeHmVl
NPktuBH/aJ5V+rrBCJzklTIr9djpJ+H4TUI7QJpb0CdC5a1n+5nT8XA6qXTFQ+TN+tpg25ewnXR5
tP+AoABMMRl27Al1qCqKoZpxx/+WgDbOpsi6ddg+2ovBunbd9PJnfZifPfrJ4MS19w3h4TsCkfzY
Sbpc7u9s4nS0F7+S/v78wKA0EBO9ZPjJ1EW5NOn3HXbMZb14boxRPKg5IcSrcLlY+A9W0jUIbmGd
HCkFP962v6u5jpKngb80LZ2aBBfOrim45GdOWlP4DyIh1paB1jw4XsBGpnumHHHJ4bx9Z56gNbph
DJtlrr/EebTYCFWr67NzUG0Ne+egavTwCITCAfJ8vilPf487h/iY5MNBKWxibDVcUIKR4p+zRk2I
ZQgiLP/Jca83UEoTE+1bc9PoXJKGl57jOdTCqxzRABHs2pg2Gv0GZwGFfMdfN9omkpwIq5I04QrY
vJJI7t4I5lKi/OfESqslu9MFBE6axdyjsGvEysv6TSzptXCZYt6oH6VXyelXzRK+TQ/8z9mdNP17
5w+CrYldU5qz/tnvmRJtwqyG7fXc5xovSpVyvtd/Nvm7Ri5jnQsk0fdx3y8ZV1r4MHiLgJy2CoJN
YNr1bTr8UEHBoTTKPoV/HvLlJtXPaffDkGRiEGKSfol+/QEvH9p3RUhMALyAs4sWmAmraXMcivYk
ZDDHXE5OZ0lJ6OYuDc8W9WPNMByJ66mXadaG2bo5Rs3UuXQ7SuPQ++9uFR/daDGqIWD6okWYwKqX
/uIu36rjbX9cSCCMDulEJNNfGtmoQNEfKAd3OO8u0E5eKlLBWiUnn9NMRyi7TUnBz0IFC1jvzAoX
ekATK0bPC0yNCKV5PnOzxyuWe3w2f84jhQ4Cr4fimIGkNM8DJ+7LkTElZIpa3/8+r6WU8jBjkJl0
svx6vPBRnVvu4uRskocc01FfLx8vJSh+E9P5QnMKsCMqe6/vdUQyjH09vVa0CS6OPXfakgbIkQpN
xnU2ywPCzovNyAToSlWqWGaayROT5uAWriWqzZxof3SU9ZLZ4KeYHfJQh3+lbky204NZq0ObcV1l
Wz+XlMXVdFz1qIj9GlHL8wGierTIa5uSxZ+Y7/d0dad9SZsMaNc+0oCj4cYmop+7LPPCK3UfI8py
ZLw6WZkia3Q9hhJy74S7zGyR6UcLDcX/vHAPnEnfVqfUbaLiBIZHpXwwX771nLNKCcIzDFdNqB1P
3NpOjdLG1eVenP3tlbWulwUjMF5cwaqZYe1RwqnPz/VfiCoLthpX02sSSozAlmPEpOhJf/ekxoR8
qhfUi3BMyvxoje22NVIrbXSF+QYLqM9Yf9KZwcj9RbCK2vWJHN3eZUtt2duUs413ArHIYmnOKaeC
2VBYCPkv/oxnuh4ut0PGcd9FzDgHtFhb6Z216S4xbbA9sdYSNVFT1whiSwLxm78NiTj+KqcbO+xr
aZ9mO1YwZNSzJAsXbMJFNxRa+pLUyUHYnPuFGaxNV6XjgAkLGotT3SEHeExe+tN2bPkuGk6NPPaG
tzZTHVn8yoSZsN6zDRs7uZVTrZiD5jQymL4N9h/FFXJ07VnhQrgfW1mRccpDYi8mP5+bW7GDjK/s
5ZT+ZBZwJBvR7bFIrJleGtrRMcGv9hUXg3qkX+QHl7DVHhcyPiOF/vHJ2deF7TTIcIwQAd0qDjtK
PdmK+ggZJzx3eJlfcfIr4UhpZisYbnKKJkplfEL7LBINJlDcxZtpo6WsZrQrFIGQg0Dfxfh1Nn91
Qn5lz0wn9TMPW6hWsttV4FAcDmtbxuOmgxj+p4gnxKebr0/vm79SSuGRoX3/pWkOUpBYGNG2l37K
/MUuQBLExpeXav4g2F6sIYfgMFbXU6qRC+dxFPmyjNW+KsWRZ0+mPic8GqyzYEJRxbhLr/1kN/Uk
oUiwKE34t6g41BeqGjMnJgdrKxVrepzvbObEtPPxJW8jhSu1TknRe5P+vjxLOm4Z1CRZ+cfLD2MG
hAYANDnFchpo9HsNjBE0n/VOd9u6p+anC+6PXQWrkb2r1CteooiKDUBo2cpJZu5SVO64NBZ7UWW1
jMKKBANXxx76xegAFRBu/vgi8YdlRwAZsu+w5xnswJvTVbxj1QtFw9O8H+yDgD2pKUeVB6Tod+6T
H1PNGykm0BFWeLh3IL7YvicXlOZMqJV215vR1A8zJ5CpOzcaW5ZbvuNsYMTZgWY2S4YQJ6CruwVj
QjYn2+ASznkyiGe/2rHpVkwBtnamO6RO2vu59yBhz3hmpM5q9pwy4n7JoGpKUrrfm6qwCHvQtaTU
ZUidrOZv86MpnV5mLdTAf9wGqyDetBUwZvSuGUk6ejWGRGvwsKwFW86dcH6ntrlA1vosnHJUaekU
a2zVsr0eZG7ST1vDi1N0Wbzg/YSbz9BlKFQVTQi1bzWYb/vveWWYHdqe/WKygl2SGLt+HuUZuYGs
VhgmwbvfxVj3mr70TrSPswABGcDa/ldp8g7F43/TCgpT1mnvV5XFbOQ9mcnbtvxMRQ1eoEX0PTY4
+eRRTW3LwHbyfQQtxzwM+EZAVRjnVJ5c6xnbGnwJKoWnHObBYCFfrI0twcsRTskbN/DEj1lPj8oM
7moc5+hNP2LVQKx+hERIahUm021BGzlzJT4wclOcm6t4RdrzRWDvjGXRQuPI2h/y0eQEgkPOwk42
OOz3RDblvrHiuZxQG+zB2zG/4SRn+bZt/HxcF6y4S/WDTuV52ZZdZRjxVMiH7QU1zWrOpYssHJ/6
JbBNC9Rwomr2MepUPb0GKGNhzy0qyT79sLYxXYSUj4ljwW4yvrButi8EdZTCbSRW8ZHhNMty1MyI
pPf4ixfsouArOMM/IqpY2j/hcJHZsfmkS9D7CaOf9EP1PP87TowDZepTxIacUI1cBWogw9GIRQsb
yqqsiCNBngn/sVl7GHfKBJMiqEuvHyltZj4aiuYnUGNEv2/q39QXAOXm9KwfoTtSAN62+oPqmJT7
spH+pNFyuq7Uk8WpkvRcBPbO5rfLwRLNVfcxtaHMeD92e+lwpwBT/AX/k7C7g0jKruT5bp2gleXR
jUy2Mfv7RG2Seml8/EsUKMlHMliNIq10bqlmksTMMxnawA8gJ9CYWxFhySk0nqm+yoUteoPHUsQ5
QqghjQzG13VtTHefgsoPfDHTModX7pXGFvobkfdc0eKLxf446dmvMxZ65sHSNxiOZP32jpszNCaE
e1eHwYbEHCWQAYqiI1Z+bSWAeyd3IJTA67xnpQLxattBlBQwFYjMKr9CU4yrBmF/EjmBJ1W2kzbG
RaQer6CYjtI7yceRNH1wBMF7GHjdCDGUAH6552DjwUBp+NtQsbB6Et3GViSPkCASj2K0W/YahBQl
brrW2c7PLmKhla5zCKRK9eOCN3QPpMg5iEv8778+EWMGpP3zu85Ma7iLxb5CpwUxP45kzFWUkgM7
TJ8aJYrUth+guC4PZhdgfOmdFhNlIQRv85T93akQkWHY0xOtlwxdw9La1Da8/MSNG9OEdfQNnuIM
W9+/RA90i3QCyNg4G4h5UOyR8fd/GQ3wROEpX3HGgusBouXCZugtDZeAAR2D7xzZZmDbEQBqe1dE
kYzOMxUc0+PEyJlSu8bCB+t6s0u4zOUSh7TNZKhCdr25CP2FWPY6gpUxCeWeWWwHsuSkwiB5NOuY
9SdqWHG24dHrIDs3G+P/gDZPElS1hYygJoKRGA3Ecpb0J5G8ay4DO+GVwhCcGBV09/i5ZtXtwG6L
WTEnuUXvvsWmsoHR6G3ujdcYo+BftKi5WYYWUZoG9lCyemRdz5rkCojfbUNks5b7zRGsTV4TssTJ
peTu1K2HULpAJxfezOdGFTSAaIQewyOwO9Uo0fvx+DUeevR8RCSML616XzJAauf8r8ohFln9b104
PRChItVJ4ptxkPwnYh8J0cMWgTXWV1k2oG3eC0HIx01EooabwZ/LOJii9OYi8Wjf7SMR+0rSejq3
pL/VyyKek7+/j5gUd59vO+6lSw3n4b+xarAhdk6cF5u/QFexSFcAek48kpClvDoQDehWyf8qJv8O
219kmmlSo7A/p1nPmsGe/V2SHLufigULw0bNE4LXeFYBKRxzndSFp0vK18Kl3qaHib3X7X87lI7N
VFudTe412tYI3z7XmEddRd1blD1Au4JfQRfYjQPJE97DF2rwM7tFA+ukqVM6pE8WDViPrLEhAoHZ
JZsdLcb0pCRWwkbLjkDlARZCwq6ae7Uj4boJN0B/rGOhK12Uhzrb1RNqwb2dHeEd9f+xRvGYLYnW
s9gpU9vDldrjtIRM8RXnATXJgHhPTYBMe+jPbiiRlu6wKvDDrhYo+e+wFlbWj2bcy+mjexfgtRSX
YbNHbCzzVe+Vdf/xA73osj8Ao38IzCqNUsBtLe359SP8Ef453N0JHUYFIjRIOBj05Po6Zz+yG0Be
lqAA+xNC0FBz69woN7DSueCnoF9WBFaoVE921WNmgeAHCN77GQKPESpGfIlMZHk/ApPezevtReDV
pLOwlDTysZCGuY2T1ikL3q1zRdatPC2aQ4FXhkpocv7MMw72exTlkTrYgR/Mln/rFGdxeFCSWPqi
MoDTMKTJI3tCNHAcu7BsqkyA/lZE136+t4DiiXvAHJIwfg5DWA/6SbAsiKWDlGhyCP2w8oLXsOn/
GJefaeM9mzYSYQdZ8otzGZcZBwqebhczGx1/LS8rlJI/t2BZWscD1huHiqsAjM2TqK5/nPyvoMOs
HBTG4tRC8Qp0F31sD7Jazvo/TxyUu1Ach6tpn/SHkYw6/XM5BFT31/jfwFrxta8XvHfiR0P427QH
l2OoovUjlr7YBsWXArpYglTmNwB6KygqsgTOir8s7EveQLDSiZiQC5SjJ0BwdTyWXUiISoAnTXYw
QbWVvwrcQA9e6GTiEdcd8ZG93iXwD1+5tJdSCTcXCJK3EptTuxAlzYX7Edb0CyLoA0Z0gELW8SmA
oqJx5mgeK0/4vw+yuSykd5dj1cUZJ85BfnKgylsrBfXDUkdpIdYt8tOMm0nj3rPrUCQIb+SvBq5N
WAVXNpU7M/tgF3lX/1q9vV+gR48aHQjDVuDiFsusOPeAxHia0ud1ucKTHkzT0l0STNSrfYnThy6M
yQsAyGTpQK6x5ytxMbe/7U73Hon/I9WZZB9arn5ub6hmWsnwE7oHBLKZSnNwT5vaIthbhew4ypzy
S0BdaRVTBaTFy84hK9ueHk+n2pzBmFaf8p8eat/WXch7Eibh6UwbzhnmBKSRzYMJDe7P+0ody+Zg
mIF0IH9FeZjZlKOgM2A4slfHQSAEteAJ4GycFHCyj4KZMbvTAHefY7iG7FCoYwYSTozVV0nT1lYO
x0Vq9dcYacxz1cQUnGZ5RzNSTs+QsVQDzt6lVbMadDIWJC0t0oj5Ns8GCpNnfDYrjBEywRcaAHkI
+aiprXd4q83flMbrC9uVd1HVSzVWj5dgnQLA9JDu6nWJ5KL1NWTAB7ntfzSvWZcPkPBgwtG/2kwg
Sq/L6BUAMrD9sCp2fTUCuhBhb9/GeX1SO8S8MXshC2YugPZDiSJJCVZFtd+sQ4FSeCTrfjE5k0Cg
V/eJUtLxF6KC9OfCWuadmGn/y15DkLSwApxm3Tu//BsRegsW+TeHQgCs1Isu12t8hSZVwuMSriMi
cEhJE54DbAazoVtZKCQ++73ImO6dUwCD8wssHSiRKvc9UQLhlzGcNsnub71dC7OzrVsKL7xihw4d
RemTZtg31FmE7mfPUCaxYJbajiVEQoSoYFPYGLtZnyRkyAVmDj1lm4lnZcZTBrop8lFN65UKNrQ+
b1oWmBzAuWtfxOUAXaBZN2Eav0XVxjSe5pDnoyELQIlywUO49AfjuVRSBYPrORV+m+lT4iSS9IFE
DbkbZAPgd0WYudlPC7gePXSSrOJgr1tnGerJWfmpuqsfGWS0Iy7lG3pVw4RvbVytkjF9/JlSGVm+
0caZYzaUfjqQeOIwS7XUJKFeL/1amtDTJ+qHSWAFlh2R4YwRC64lXxhNVq3Y47vlMrtP5zG56edw
iXHPqKvHP1odvd+BhaxHudw0zA3p7Aqm5jr8r+1QCij2la4v8sz+cQB7cKrU2RrJKaTCoui4zMVH
jmF4Dlbb/cgx3oI8LfpImmao10d1HqziWgERLh+KRH4O71a6cmm2Ka2tMPmjZjhqRb/rfUSVIKre
CugCKLXslJ8JFxU+Agem87YhQMSHgAgFY0KAGj1dH0/EDzJviNZpDXAVJXvX7oek3t5RhzI7cwvu
w2wJ04nZt5GOv7lIR2hlIzq/iWUHu8njnEcHNkfWRfo+aMDPdzzOc+jQwxxpPyHzRoxqV3QzAW6l
5RQ84zHfTa9wE4Te5xKiFHn8s7jD8a+EM9WXvcgxVC73afJulFx6gfcwKU5tnlBIHBzghT3TBW/8
nuVTCJZCmITX5+jhUKWVIeyDfr8SAWZ0LNyzOh/VmgcvsPaQgLwvUvszgLv9pt2Lqj3bR2igCL11
9PiMGOuRtpEBSeXXrMmIf0wsUDVwBLqDnxbWG+yokXSRDl5BPF+9bLqmlOADsD1x3lm2MbJzK72x
JfD+RZiLXsVpQuv48kU9HmhA9fkWYZwLkzbB6VbeBq91Lzj3jEjMOVqR7p/TSn8JCHaGdpV6sAl6
Ia6NjR0FJN0PLvIOxU8OCMJyj5C1xaFOaaxO7aSxHJBw5VjXOgc2rPEQ4ufnJD9Yyzv2XlcZ920h
hDTIYE6TjeYQjhYqLF+JeOpbuYjexOS1oAEwjcbG79A2Kvz/DE0l5I53G3xYIDPVSqVba9Mj4N+4
2wDBXweD0KQZ2VRU5fj+h6oALRlKA6R8eBHfr0scr70BpDJwJ5DRJVRNC58JGDLRsJaIVI+fxQzW
CR+c6xIc1sPEqy1tjcQPYlCiphs5S8Syox1qeKYWnqXRI6SFiC5tJqxjcRcW1oMeVvoUXkaVW849
DjLbyE4CaPGMfrRkyKAgFR8mq4ADlyScO0Y6jCPBq/lTmcXyMlxyOrEUWH94Bg0u65JliBeDP+yt
T3eVybTbzSuvsdO87d6iv6f3m+M1CITDeuaLs94gz5FSuDEZMh0BOaoNpPIQ1d7VoIfrfbWjksYG
maZcEwr79FvlzY387LB8vJrCdI/ghbACQG555utYf2WX0OT9eixrTDGBvHgBMI5nrrwpXDWFNGmz
BRcnZGtvJzhd0pgp4p3VtTOw6Nn3i+u+GvjiRmSirnikVf5fui1sFj0NlSaw4IoDAvt5eCmwFWrT
2TU7PU4e/td8mvjg+XiPkkoBkudm+ltI+PxoHUI90M7FsydnrV/SHkOehofIpbAxwHZ0LvljqXZB
OoY2iJJQ8lOdEocAXado1nLvWOnFteDWIAktz0hgiasBzFSCYSCTKcgSiwsgDzDeQcm/3gSf+qG7
KeXumioLnhNA1JQVUjIXp822rXnh23myfliTnP/BDVehlo2WKfjpDVuoEfZJRjd7cHjEkOEbrXr4
vm/6aLRn4qtr6JNwKXFr7egpqi6o0UW52bu8+yhTwp3ywsPvMP85qbgLUTUpX2IXfHBP7A9qDY3T
s3fkKyDnRR7OVMipDGYEEVIgwcOZT+4XyBdTqRlUPppmWQ2FOOieY/9Yx9QT2Eo2w4kFmoGuYAsq
eQZbGQzSdZsHPMp2p/C3Bs7UzS/yZEOGR1hU0SbJvrXWEABFN8AzrY5MBlOQ3JYqk/lgHM6NsIHW
lXagtCwAP+XQ2G2cjBQgiM5gL5grrrAi6e4peJHkp4IwZ+dBezygo9Wt/XIYQfbWf0X6KSpocLr1
yxubbTIb4p/yHZTwmbwRMC0eOPsCb12C6z++unbyLXZc2oesS+Oe03gsFVFy2+YHXlNrGjVaKvAH
ALEgEOA18lmYt8/Ct5+ofYYeCFoqmyOZwjB019Rv8+2YG7Zhca8oKlk6QlakySyUV7DJVT51OlTf
KQzLXOC2vNgpG0msQLv6KIAPBUZThqa4aKDax+AVWSN65Huo131MujrKqPn06K++zNgQMi3nzqFf
ikI8L19+vBO3PAGbgd7vBu9TqZM3tV+dh1orNYcJCK1XFsj6EnWBxuSKXAGbpKl5aej8Dl+KfBvu
i7Qp283UHN1ILaaZH2bxQQznKyQTA2xwvksOf5Fr8nS6kjtR/JZZ76TfkApCJmV1GG/nBfophEXB
RWqx4cUU50ZzwNqjw7HP7iox+65M0FsptIcr4B7NzdeOV1XPHXSzxwmSUXeW/zTH1/tennpnCXtw
0bD5Ynm76MTXsy1j+yZFSXCqUM8SBraOixTpF02/upCkZ0mtNkPuyMlgXtaSvFiAutoFJrVDm9Vk
oC++6p7dXVpbOH/17ad9W5sXC9m2Q1le/9R8Zp7QfWmFJMRUo4R+pdh8yGHTdYO1Z+AtCPTB4iyu
UjA6ewLQgFFNdtB52DSIQRRSTppGDR87HdtHW+8bxQOqBYewFYSaVoIOsJE3TtviIoqaLyIy/BN9
JUOHeFopZTDhEtotm3UgT3IYg1r680PysuPaJ2hLxgaIhSXtRI3PI+f1kxXQMMe9n1NbhJe0g2GN
OosqIz3tCpoMBCWDfaIXKggtF1y6+e461K4pUxmEgMoj9ODkIUU3NJAavKm1N3kpDE9Cpe8TNaQF
Ctz0wORn3VqWc1U61W03/ji9P+KqmqPuGPGxO02aCBYJZPJ7XgNxCB3JaY/6H/kN2ucV41AO2f3R
mbjDyGMlhUmnIkVWd21NmIpAtYmm76iP1UvDv+axM61oudXrQM2sY98aB8gfqKP21ERHmgZdFDUM
qAD6Vj2dCXKrUuKz8QZ1evT0tUmFi7oDDj0yePTiZxvoxG5DICNRUNFVKQD2y0lqikfEYxFOhySm
VzIZh0BAFEx9YdUbpwX7dtT9SXyn5foGecJFBydX/8plHoj3juCnN3sn6/lFFcR9cvbBL3YcvNDl
YS8zeaURBfsRktCwk8WDKkwD4tvp/hKFoMnBJNcDVW32A/Y+bmqpuz1KQkmAbGcIymfobymUjUAi
mkb0pnhSci1xDhKRQZSAVlaPvsnt7zPdJvg29twotx2NhouQwnf6kK7wev62KZHO6ilU9KVmhiJs
njs/g8AjzTWRauKTLV2/FqzbeXfUT51G8l792gleKxnmygnJIkD824tdzTUFxYTVJ/lDw2KdBG20
iTNaa5OQCATPn7K/mbwv6DVhmZhW21MGqIQAzzBTKcw2A36ZOT8yeMniksZyblx4dQvD2HbBgmeq
uAFH38saqrJygc4BVrYehcInhBSL63130kkzapC+/nOTb81FjvutKDxi69CztrobGIWAeB45knN4
Mi22t9MVaDzDP/AC4NOFI/XYI/RmIAxP724yV0UcKkkyynQ6bdYK0Rah13FkWlwqaRZUL56i2xPJ
AwGWfh/Los3CSw21IrUO7m1bEViI0GohR+0hPsY48Lta3/ksSNrYy3f+x9Z4pcRafh4gh5xMM/YL
xVTt8/gvIBa4cd5XMf/4rpjnJfnBLgHdQrha+e6aO+pbbOtjrEQzKk4ChoJUXk2YD4E+u4liCjTo
tyIT7mTjqly/KInCN8VatLz4HFW8lafFdImBPMetYgSFxJRVGHF/vAZKKxO05O0RqdOAxrhvM9sM
WhKzJSyLEnfJJgoHHp5GnyH+Qcumsmddk3BKRAtGr+oh6Dk8ZwJlL16sw6c83zXHBRFhMk0m0GK2
VVg4naMR7vv/EwtRXwKPMiYukbLxntZgjsqQ5gyuWNarqt++RzkLaw5QixF257QOv65Br3okUDPA
rbfq2e8hY8FipY2v8c2S5N5cIs3qiDs7FuKfW0RmE98Cm7v4LgAYqATHKMCxnP/q97aICwD7VmCa
L6CnvgpsQIvEV9iMCCX+NON+XRM0l2VL2Z21PKa2eXJbiwRUF2xFjfTqCa+uT2juKjGP9YnU65bK
B57d95FqZR6b9umgTJIMdSyCQNxFZuaEytuCScGpPom6130Ju4aZe9DBjEDUy/Tq70dAu2yguDr2
mXKIMbu/H7xcy9L45fZXZFghiwbsc/bVcza7ZG/11SlNWDNq0EfpAqUI77CKzRdOmVPZ1mEiZ7B2
7ZdtK+IF/JGu17sq2xryYJpcQGOYCI39TfV8c72+uA9iMishjFIXV3Yo+4o/fCQqCYmu1hnb7k4L
x6/uFYScDHmpHI2e09f6mhCLqu0ogqa7bPPHIrOYx83UK5lZPs6niQHWI9OJtALaiU05RmF3USgt
777Tkl2KFgGt1sUNbE5kj8ZPyojlp1cM2p5kbwciRhP3bdvD5ZEbeN/xCl1mzGRJ04+RmXgmDTDQ
R4yUqk2rgyi9uM5LF4qzMHaILbJGe81aYqdlNNdp80ferbEIFdktgCu7Q2XDK7/vQey7ttCqB1Tz
uWrzmOrBWjIX3uRXY05XwNGP0DNLnuad6xiB1MeVdlD9O345p017mvzoksIoPmJPNswThOSdmiQs
Z2GQlEld5mqEZCFdL21FOEmNE4LH7CUdCiDR1PpiMnJGQ+almpUkNtEX4vHz/yHSf8m41zAvp/wK
GPzVO8wd6a2CWp1gyf7rZzz34yIXl+mThSVkrQx6epICmRXytNEOpZTC32EGfA33yvfyPLOM1wMo
Hg0rv9z33kKN+BJ57aev2tINSi//SPkda11LWUomz+dOpccsUCtpavNAqFX4vJtBk99Tb88HsNaR
QCLE6Kwa6BQX2bkjS9crLjgbIrPWEtHT1FQhk9P6ca1l7q5XRJLpkFCMskIYaI2AC9R9KkNAGR8r
Q3gAIRRIxEfN7GUTAmRyv5cSpe768N3fhlDRU/QV9I3PEepxgxNTKW0tU98IdiVJ+CFO5b97nJ1H
Yne7lEB5Lh/vtJmP01gTVAvgHITQfos6ukEJEiWGa6GF2TAtCTFGVF0e4SL+JA6oH+aC4K/Txelu
65tZvdUZF3pSDDGif/96JrzivK942aO5B/hZ3nd7CrZNF/+r+AFbqQ8i3IeB+xzmU+IxvfdyUJ3W
AfGNwOAGTj/YipbQcUiWye3ubuMozmXr0NKxdW6DSiBCYu45niWnqmDsO73jlTHtVBXgLbSRMlpe
8eCKMgw/zDjLZhBJQBYk5U9lg6PVuNvckB5fAYcbd2TlpeaGgSkGx187Uit1fHNXf76y6/Sz8P6f
WdDWrVSqcJdxKr4fpwqBKf4eoeXVoHpf81/HO7rmpOuj5V3aMAupeLQvjz/97cBdNMOJ8k49qjuq
Ij5nwKEsvwvu/G3IoxnqgvjkzquoGqv9jAT9LorVn73k89nUbBtCPTdZb/WUGZyr9mXPtrmJ6Ln1
mI/RGTZ2Gfhw6tiqOSfmoh9sq4m6GVyFPMF4IBbABdMRioE0NCbMTSos54hQtsFssHCuS+YZlp0t
3qDViZKOVgxa0l7+eo9oFNcSFIOLJ2zNDQ+1ywnULOT05v7hGQ5YJW+aKuD9paffFP7FFYYWNDwA
qTNW4Fl3rSOzfbMaXii0lsFSchpzp+ZYC9KJ1fbscVcmkljFLCziOe7wnuju+F7lHgJWezA7Vgm+
ZUpemRILgF8nWsxNPMjIqJMrdhzU4P5KdgPlwcyuP9ZoVMSshh17B8cHplTlZVp+0EsW/BhpTTTJ
hXZhkvuUeeD27TT3ycWXS021eN58RByp+BSEbiK7uNbl3fGtO8pleq5tB4NaLCO24VC1RTfL5k4C
V/OiCbfXdY/eUboZusQRzJ0iFTcSpCI2CtIt/bEx0Sf0DnmyYcKUbJBjxXadFj1YT+6xs/9Wiogz
qh8UZ7UA7tszpVbCt2eL7mB6cv78JacUK983eFaR7zM1TVeSRdcZaXVguyR8SVB6Fy/YFrc9mImH
t2YnvaLfU3I+Kc3litz5XzSwieknfOjU+rkHQ9CJ4cdvOy60z0mhHG0ChfyGhqCs7IyV8KNevlA3
O6fWBmMcr6OVvgjlQJiU1Aq40I+jz8FoaNVmnf3VU5R+6Z2mF3VQBSVf6nDzrWQvQyLtGh3W+u1n
sZHoHadkmJPnlQHsXZGxucsbnX1z9bxOozaz6L05Sr0NSzxwto7uoJo8IM5tH0/LqKVGRpev1o4G
LIsYXfShIodNIr4SbjErOEQ5sQsY8iRu5QPQYvnawkVzs/wM2G40Wl4c9yXaNgH9j3ALes2MC0K1
U2qRUs+jYMW81HduZ97QD/Y25TeI8TQtowM4b3Z/dF6diCX64O/DWL2M2EOWunjru0wnoos592WB
AhNzf5h/k1pV2z/2oy5rEsHdXeFZSrhq7aqlv3uhsQaQ9+p11/nJoyRYoutEWG+budq2CIPbFOo4
M1WQgETjpRbSflvwEh/gjLMeba27MuwWcNxXCi4b3qBGAm/s+Op/ynSUyYfSt04beFvoSNPV2+OM
bpC5iJyVTKaEXIXsDPlqjN6bQxaqm5E36CMt2hUoOP7FPwThSmTpNUrB+EUvlPCsDNREDCF9AQwi
f2McLC+LotXxcSpqlOkpTwGHkNooDWdJebuNx9Z0Z6Gx8bt5dddAs0MgED6wdOe5xM2tBdvyKvQ5
HyBjuGdxI4TkLB7ByOPMxuge74FzgOxSzpQsq2UDEKvi9xhx6yEjom5QMTG8Gm+6hcpuAk2qYjk/
8XNkSQWAM4s+q6zLad0Rk1NlBWaFrnb+dynLPEl2cRReqA1T6JnNUQtOw1XhHsVPaTNWIRI7Z0QR
lODEelyZC6ilsz5CvJpPo83QcwUMsf8t8fjY/nmh22VGxZeDQBExCOLXGPWfUzZm3FgroHimjpsC
Rew/g++i4WflvOg0B3SqjIgz6Tmyn/8MJaht5z9uMwIhPLUq5BVUmOvKqKarWaWX1SMYtc2wg2lx
gd5gNM2M7YI/nJeKT7Dexma2A4MxcuPBBXUg7RC3I0uPRjpMw0BLNGELZtSUB0QaMNHFTEVhVc6v
AQn9dDU7DWBnu8sCw8VoTqs7VGfragA0qKqHYZlFRK3pr46d8hqHP+OFMXjQBS7cBgbTpeW18fyQ
mpCyFz2pax0ana2Wnfp1mJzKgUB4V0YjlEgFNQt1fV6EC3p3rXJUF4pXwTZHs3q5Aw76urV/Nooj
zNjmd1tYwgyGqx+k4SdSoLcB/mAth6p9dUx5baJD6qK0cvb5t8UMSgxTLGr/nT+/lJE7VR5C73xG
kbrGDP6OHTCzQBtuANfzV/HKOQKlciFZeSgDnp0CtHqBkYug6/Z4NG6lhWjDIN3Vlt91m/sJl7p6
BlABOY1kif7St4jRW8BrlzNUG/fhGyTi03X1QlTYNPL6kuHUYNm0aFVMxf2KcmGx32bpOB7LGZPc
+dJImKSjB01iJp4Nau7bDYDp+QclfnkorZ5VILIHTV7oWyB75FnjNen/WwFErgqAp7PPpAYSCMhs
YjIR5j3VYk6bwMd+Pui5uSZRVYSdko3K46tJtBqQa5KhxF9xN8ijFJ6SZYaNBIdaH3I6p2aSLkMy
bpkXytqWDNgAzmi0XiCOjpXu2qwZLZg8iBS6cPwYWA3jdUsZtiqReb+xIASU1rqyiCbXaV3g3iAV
SRULTY02Z6LMl8I3MKfeRo7NWuK2FvqwwioS0vMpDVdPYxOoFDMKqbJ1So3j3z1NRodCHfNRNb8F
+CK823wSJm1mF3bonwVgYzz6/b50bGk1/yyLW70XJ+J1nl0fCRFYBy9x1fPG6z87tFf/EpxAVbRn
jbva8FVupq5YLkoXKvW4gnNcFl1mzk4zEyF1FH17o+d3d6/JjtynY6KfX5NgTPXu3ZUaOK64mRG0
XdJw1jDxkiMEYg6gw2aDhwwfmcbQO7M2IcabWCl42Upq2jyyy1ovXCvg2f+BHYx/du3uulXNvu1L
el0brp7GQge+llGEklQOhmgD450ocGU/F9kLb/3NQPXjPFzIaU8W6PMWPq5HqGhxL6Sd2TZjJvmA
TgeFlGWAczxzZj6vKi/mN9LzwirvFNzOT2Ffxod2mfY2GoKoYRlbEuQhGsI++c031LP8RIzY1g56
T+P8fkUDXEvf52gzLxNz5FncJ9G615rKfCgLAuk37Xo+2DxzEMAF4tYoPQQGOxUw9vVmLC0j6TNq
7Wv9la8WKTe+VhD21rzLv+l44s7EH5m5Eff6jquCchlgbitGryEMA8BIi75/IuflYFccopmN61bb
Kx48SkWGmnRdvo6Tz5XkLEW83piCPjf+ggUO6jYcae6/QqSmB6PEfyIDtVlRW0ylj0ETCbz7Rg0Q
wD/A8jS4zx2PNacjvZwiH/hpjuZbb6A/p3U1sPpfqQWLagmmKbGuCQxjZcga5MFJnMgzLpvsdL0F
1KEw2Fg4IuE+aaYhJPJ5Xj0cnAo0Qzr3ktuI3EVwZ5vsrtETA96FPRbY2FGkKjYhbgxjovMNpqyN
+jNbXihcU91O++4PyB/W8ZNLRSOoBJp9kk0G4lmw22wFjwcHo81wFBQe7MUp1gYJ7sMW8EzLBeyp
ab4E8AD0puRFjNw04AtcwmginHtCNcnsofpKK8aQa0xrpqeNFscpnit5kdzuV1/BiS5/cnztrxt8
p37kwySiDFkvx6tL9oLnlwB40895y9Fq9rBKLLH3ppgozmm1XeREK1nLwmEAC+LAeoPZWFfT/770
oFkJaKXUUexPMZb3sCenHOUXoD58N2NAtWkVke0Glx5tYpycWtzj349m8x3k6P9sIJ53h9WWwUPh
DlTqchvcIcThh6ZPq+L9QSYwQ6oWuHMXxYTYli7sXkGcQS5od9/TqdhrYf8w+KR7NndVv7/3STLV
QM9tDHfkXR41JnZfFa1URcP5S5T1LI+NW6uhtPOy3SA69UJ4xN5FCmM3Ob7ugQrSsC9+B4ZAcs5j
jcA5JecZfOYkbrdYWjxp0gt1SYUd/OPxFTJwStwMm7umLG8zO7mPZH0ujIY3XLcx1yHe99A91rTn
PkKEWLTnrOPvH8T6vUvPFMqf23LZxgfT5wDx3bDxmqIYctiDygJoC8AiIJ5OnOmned0sF0rX1GzL
ZVZU4s5HyftKPGP/r3cc+83PiSbwCcNizXENxWnK/6zt+BDvKuh6MzeSgowMGSOpPVIvefHuZDhO
q11IQCIzT+5xVsn5chLorpzaDx2ZsaBKbunds9ia0YpbriJX/sda2rj8C8GC8v1DRlw3fR4IFdIk
0fRiYPtqFirwrTI9Blsl6/0u4B0a+Ua8lCAHm7hxqIQKDXvl+ewXLSKH0YZSAX+CK+5k4Y9uZ9jF
b6STvd4Hbz9/HrfrCI0q/sIXTyB/Scd04LTpy2QlGphQbQvcux7cuyAN6SjgUEFslZXxdri+6X3e
maR4Yow074V9G4K5k4VTJWs7iF+efKtFO00xRos/cC3XcRwwl5FuUZpWEduS6xjJgexLT043Rxps
ZqEm0bSByfnWQgCOKTYVxsTHAYFPI1RlyhMSef1k6klzC/iciMoPk20y1Y7E+U6UmptCN7Y5ZYFO
BCVYCXglHP4gFJdydyentqZ+YtViZ7XTbtwlqB7SHjMdA32dGFjdm2ZnpKR2nugGqe0l5l/S+MaH
qbSEJIYiaQ2QJ80X1tdVwLCciu5VWKt4QfltlY5mnWbBqlTKkg+0buBSdMv3iyNzvNAkyFngvibv
H1Lraf/8MKHhgKG6BzlvCw++VGjp3DFk4NBn0+LT9T111lmHLneJ1qqoT4xtLJtXGNehwZXzklB9
W6n3m7cH2NUXncUNPMMaU+tGiAo5RuOsnTVXpIWXApq44obZnnoxpXfGuN+yGN8KSRKdVQ/m3XOu
Magrpv9bMgA3SEVwGtnfDq+UOktFedBV5Z/4e5QDeHnyX9uri/06nD+RK6CySc7U0M0b4aS6cq9n
RPApx/kFn/fI5HKnTQmG3GYKHe096CtfXWn588HykTQFaW61go8IaaBxjAaXSqxO1FiYQzUv8wY3
BbfjmQEHHOhdK03qLV1lvbnT23hVYixtPP7cAmfYLRKxaRXhO7YqyiObg0B6PK6TYcGiqtZAJ8kr
tGEqr41jGbM85DltxrjPtlKQR0ZYzQmSiIbVKOYtrRapBHMmRnSk1Uclh3cswj96KzbrnSSd2IOf
ClZslpqmGlaOaGOjOu7FJuBjH18qP88nP9rXKea+CT6oD6yacv2ebPc8Dfi7Rwgj7ZLPwdmCLw0c
D775ucbS8rpqZZIMYqxTj+qgMrRX+vP+ij11g5hhetKB/zSY3kf/f2jGfp7hEtAr+r8uG6QKROYH
fPovRNhSiZ4C/w+Wrx0KD3XSa7exyA88wDNEWrIC0VCEpF4nMmFpWf/7TlMzO+izdx6Yy+uwxpwW
stnvozsio6U8jehl9jqsesnY2ZBQFhpS3Z1mwabTAMNMXjZb+r0I4AT1FmY3mmlG8FteHaK3mrld
8vif5Ll3RdMql7YtsevoQMlbtnpbnJ/L5PnoGd4ysfkVMaL0HNrrJbaEbB+ohlgePYr8B4S/WFPH
bMf9FzDbueyxOInRBqEzuKsAA+P6vnNeu8pVHmLqIayPeHIPYdrQN33XMaQ0781rI2qAJUYWYwVS
EyF9tMVO2KXpuKJZuXUkGpnAtDHHe8UlVJ967A8NsrIxKcMZnTeBTO+UrT79IF13wO4Dhs3/WLld
ZzUkhCadTgWSzP5vAbGEICl756FWxXj1G3ASpHZwf4spT8Genpq/WAXdGd/tlwbhPeimNT6JO2Gh
eg6lt7cjvuPuSsm9pieVx3Jxf/Sf2YvKwe9xVn3CArPXOn6qSZ9WzPYgWXu3FEjlkqxyTZaEvdkf
zQboGPNgYzuMFALKeP6qLa9VU8sMAUheMod1Y57/kTwf9rmz3Eg2toNyljeVAmNBFX7JIhcnZWZE
c81jwc/Z46bLTcxGjIylBBuHjwJqsPqYn5wvYnNQui/OiAVmSTWEUTdTgNyCWt7QFIuXYKJl3dPw
yJW353XmNzjM1s3xHVPZuHaMq8TvNc6UDzFCzaqkmVQGqqnp1JYoz/9Q2JsS2lguvzNy8IVJqjQc
WSulLT9v1ya0Yh4LXYAik/6ykJD7NgRFKObkytXuuky3zm2wPKBJ9TasHxqoGB/gARqYg3QVd5hp
9f92xndKvUNbzeIjK5cBdCeKWXNedS1JM0n0lnycZ2s0mUMwIOnargmsEDbt1YUeA/aZ7AQOXElF
SCfaELV0Oghr3kZt3QLi2EelTx5N7Zp6nKUcYQb82VD9tWDsVJNy2Wnw1kIx+wmCQnAK3WT+x8tq
3d0vHMWjOpIrkss37lGESICD7EMgKe22sUPjX9wHybLr/SB7w+4JpXgtZeLifn0tI73miITDMEjp
mf3aRcEHnDV2tvgVy5d8TDUngapu7mcAQjnlMnvWJA1oN98c2enxF/iH0j/GfQv01mFeadn/sEWp
Ba/Ww/w9CNFYiEQ95EMqK6ByW1kXD8Iv6Fzn239hNCbNwN28OlktUkPdaQSwtJtL/oLBuuxkA6Mt
1SbTlfJr9UYh9D0nzR2JSp02nRbfO6NTjNDnp3/nd1p87BEuPG1w09SHbOOy4YFa78esfclmTv1q
cXFbSCY1pdQVLuymvOnDsftxuBX7/Aux1At73vlwJgV9CzU7Q0VoBPAAWeET9G/zC9hydJkZLJhB
BdMs60pHOAWCQIB5czyT7jYNEYMbOJxmacs00QibDYxXMAv32tBf6fWfPyqY8WUBDU8RAluFKs4+
Y2dGhVBuFAldazuk00WNNJm4+lzBXigJwZV3hvcSWkhWT8nUvhEcj3YR7SlnABuixyBjK/qCiNLv
cYdqfwQur5be2e4D1ofo6MiQu1bPukf8bGJEU3LC6SZdJ5drwjddaUsEshP6tkyK2qh6ZM+9GUTn
aeo5jCdUR22oYRFc4NG8wtdxo/mgG5MORZ5ODa2ryZKaR/xwtcYDK/MqtpblSSCqRLMhYPJHwL0+
Yl2+nKKsLchH3pXZ6dNdkmmJlQu47SPJ/ExQFR+gmDC5H69EH46b782W4PyxBLAdFIjySQtX/C+6
LQF0zKLRs0X/4SzNWZhHgaDhMnSWAe+A/b3AOgXWu9Y7gNKv//H+QSu6rDy8yxrg89nFAtBHzvEj
z2mpTFChifTeAYYSAIm/QFXVNlayBCv9Qx8t2IFYCneh7LRPeV8m5OZPO+ogZ846b9JI+5f6MzEO
8PeFSwJUhsDAWS2ioL8+9SOxvVhDMSgntk45dN3ome6azsou9EqEARVUXXbE6o+H2fy70v6ZO4cu
I3sI/dowVIyhZdptZiGUMnPH8bQpEpBCmK0ue08M69gYxWQYluPlHb2xAWTLgpnIM6r/pMv7ujo2
SXJEQmYlVxw0t5IibwBrsaMLekfGdphSvgaFrEKkcEI/OG2EMVRxJ8ECjgIjHl80Cl0E2bIx8JN6
r+4Or+A2Fk8BbrVM3OF6QjGFF91crH4MJagmL+0S7FjUl+A1WJYk9QD/qg5WJkmuLmaxqLzRrjXq
0CKDPTx7Bd7XSkIl/YHAYVYNCZP9FOVHAJs8zp8vywNwnq1XUkS95+5B0EyDnISJBtvZMc/c6PHN
aGlLI1EwV8Wl/T5rkhe0Nu75tM8A/lnHW5JAZ0vTr44ymKtvuDXPdEwhSADsHI0yBb+AVL7z8eeo
TV5ohEKQB4srO+R0USn3HLR7J48AeQ7l9HF0SqDHFlkpT59R3VD79YBYTCw3uuYBnIB0j1I35TyD
XHP9ZC5ivRy50au9rqyxYn79cvWiiPuTlcyrCBqLWhhdPJrWIwO4kLfDdX59EcX+uOUgXf76HX+Z
ejUUMDj7nh7mQnaxvIrpOZi7KoRoqJutGIWRHZKTh7gtNsP8qV14tlMMdLaas0aIRZh1250Nw+oJ
vBwwvNISbLn0yHDuxDAcroJojUQRvVmgIwgdpX5tmSfo0qj9vjnHnmDjIPmW/yzC3YTsLiZDpR5E
gLvXOpSSE4MhDUOGfZNnT984G6VUQ1WAW4PgyGCvZbvELYVeWa0yqvEU55gIYSlcHyr/OV0ds/zU
JzNfOqctr7wxXuzXJYTuGI20ntfT2WuulE5+BA0qETA5Jzz8QggAsRSoyjQZ6HQ+IfgnbzBqcYRc
lnTTRik4xaM1Q/YvIVH8+KgKv1feSHg5RmZY6m4yeP9xuqujymE44BicQB9U8mHCfeJ9oEwRMqgn
mw8MCk7yz2oPoP2k2egbd0kUGY35WsMHOfLlBh0s5eXA9USuJALRr/iWwU1qLql3DG2LgOQDG8L8
EKdo6yJ6o4kHJ1v3Py3Ek6qV3kEyWzk1Nm/5fDL+jVBuoXeu3yoQT3cIFz08yjYTSjgCdhSKEjWK
IszTgxUeZ7LCBt7KJAwjnpadBm/lsyCPjrpFJghsn6RJI7BlTDOvuZECq8kRomToWv6nRQVzGEFn
XsQsegH60C60CFlSI08i9ddCplQvUIkxuz3b+uFWl5VA3HE2KYbQonzcWmpuBSS3Y/ojcE5h2ufh
fNiSC9c8qjYgSGaJOH0Q/5j+beS/v1A64zy8YXFvu6uEJATM6qJoE45DUtxJMLQlZrT7cxiTOLnQ
QoGYlU+XzXugqT8fT8OIA+dl8h/7ED1rrDwH83WJMZTVDL2240jmu8/hhN74pyv4Vw3IGpjGggsT
scpjW093fBQo42bL4TG3wuCFBAVoUd9ooJnW0uzKBmlUkcxSCfKktdnZXzQNqlxQHe5JURbo7UGo
pyRbGeKaFWcoy6gC0qvh0FkNzwlvdhbPT4dqD07eW2/Pl4KkqFVagd8ncTt1051sbn6vBDyXUE0h
F1rkKvwVpz9oAMiP/Mfm34M7USQ766LKOrGeZBVAnZsEjPpWGaV0CPp+80/a233AGLrKwv9SX+cp
h7Ww5yBKMh3O/Fv96KdRZnouLNk+B2+mei3DQ/9s07LP+7sdfW0KsN8Gn/gaDI0ImV10ai0rZ9E6
mv+ELpb2PpGM4RqzFkmQxnPNLOMZBtyilcPgAncJ6fwXi6Is31lkv46eAu/Yvmg9415nIlfM471n
NsAS8MkgLXS2C5Ne9BC4hB9Vvi+F7wJ73ugtx4GQht1QbrLbcRKzs1f0oD8muwo4SakKImB6jKXU
JUyamsdxAo8yZEySbE1Jog4kfLUQDXuUnLBdk9XkoJSM2J24BRlOw8m395vPxBTZwpaA5JK2qTe5
H1XAbv88Ese4kASmCwIT1mj1nFhyQKszbkiKhf8B7b3qGMEXoHypF7AGtHHrBZ/lho406kHYHrbI
EkcT1mBJ2mXQKZX0JA1PnF+kVPVI1RZITEW04w/znALn2Byr67RXE4gon6m+q31ipsF+mxlS1jB5
PcYYcWvPqWo2AyLj3qZP3WS0EGWGDTJKFSRlysS1lZpRMJNABK70BMD/eseWBMZr38Om7ZqzdB5O
pvuM1akHk93N7WdU8jrm+sRH6Mf7vqhHiP03FO7lFdPXcIw0WYtydvYHk4iCEYbEW1D2cKpOz2zW
8D0iwtVqY20WaFtDhMu5YHCbhxWsQemNFOm3x3TYPLbUxdfc+elKXu958sRgmxwvpZ3smwCXtfji
51xv4Wy/gFs5MHnfN542RKrzFcUbXjEeyK5974bV/Z19qRVavrxohD2GLwvNCcdO13B/TJrdPodY
FnnIrSF6dOJPg/Eg7nwM8fQQZHd7C51AXGZ9JtaXhh3UTBVddzTWRV/TKiNc78i2SvRRNmDmjHmr
QjPgX8K5DJGzSrG9WBBEPVC+GgkvKcX1CxHcSGGMW8rluZRiO9cf3pcPU4paUj7op3AJfvCiXhQX
4kNVFKuV/ESmIrzR4ozR0EabsfjLzDwLmgUPge5TqGwKvyrgUX4FRkxeW/G21V4PoQVnw3afmNam
wGGMF6yi2WfdCHcHdQzFAbkI6j9hAHGn81WY5AMw19kLVVOi4qLTZRreM72mvOgB3KafaHqTpMrd
uUyWlIwfxEGcwJK9E7fdN5WQHZbjvE9En8MlSO8HZ6z2VlZnzKf/++5akTUpYhoZJ1hwaWVMw4yi
MtbD9ziQRUvpmntdCSDWvRE+O92ETDpKktFvgXgMV7yGnv2oQVUJQVe2n37R+NbNUkBbUaSWj5Pb
siuRTvvDIwHLW7bDnudrhuWQxTRKaj4dNrRcfuArBDplmM+dWXu8f6OyrsPaiNMneCYxESwlZI0r
c2UFrSu5qnlbzaxI1TbGZWgBHUUvVj7AaV8utOD7RsEz+Ji3SM0YCMm/8l3tcMDl6Vc1y9ZYpBRp
osd4u6/Lr2NU4+AUVupG2VMnQobf3MXhKjqdevc1eYqXcegk6T9RpvnA5MY9nbl3dX7W9cVqVxlJ
Z6zIw4kjhSH2BJaFk/K2jG8zK7hdC1C29vdh4NRe6vi9S4VYkl+7FSp/td4zWAvmkmooYFKK8SbI
1oFZ/2ZtGw8k9YKJUhQ1vpE4dzxcU620ZIich0Hlrb2OJTbN3A7p1kh1iCrKwhWehbWm+WKQbKGD
VRpHn98iysF6wo5lNfq9aCnphlNVtK+bFdXghLd6FblAG2qtvpLfaOiz1rFTLAAgwYvHNPYMzxM4
1Ci387okAeeKoDJGlTRpO0MCFW6Rxcf+SMk0NVdPii+E4kIzyoij5bojwh4QTIMJP8zVYliuPik3
S/YW7VB8Rm5qKRKD3nXLhHmB7diDtNZihw+2o6ZNw8xL55KX4Mw3iswkqrQe6+LCuUorwBRbR8Uw
RaTDikgDf1mqwOmxQEmkokJr3Hd3KB7HQ4N5C9QnS3IgRZ7YCl4fWXvRnkPO03q59H2Ps26cf8Yf
CmgAqpPKxn0V8kFBn3BLdVGxUMEgGTrYzIK8ZeKAaSvcjS+wr59/fRvlZTzbqpFRDhY+sbcqYFxk
6Q2y4Z88RwQcSUYV8YHXGrzMdyJmAtmr+cews3KnqxiczH6PUGzh8FBEWM33FORe9RZ7gTZyrSuf
ZBpC9gqR8SdwDi8m5IPW3o6FkAPab61bKlqxSCS9mougDvZ2LmK1e37z66gFlq7Ppkh9PqO+OIWG
LJ1onMz4PbYqGWjanxC+FBodmflja7G4ZAQXJJs6j47JGrUms3PTeu2gBsf6VWzbABcJk+3WobF5
PoH8TBOfmihxHtg4oq+P0D1jxcl7r21mfrdMDkp9Peha5VHsTHmNp323URMpAnxkXxf5TK0jSTgg
bS9cIBtKoXEOM0sVHpKOcQ5UqPhZ5Uoa2npoFA9vVW+UWrwlScUIIL3QS6FA2nqaGUoJwso27X3d
sJYJ2+7RJ8rw0oaPKQX6img2xXbdZt1IXAoowtXBhqkt4llyzH+xn1AV4ULy/fr9V7QKWVAv7ZRp
E5bwgtqglObyy9kDCi606cMcs6ggDsldxKLdNwBVzvlYlatK7YvnWjKC9EpWh4A/TSp8fQ/BlWpp
6BbubE0yH8559ZAQXav7C7c+S730pMXNdKq1X5p7AuvkaafWtPIzi2DtY6RT4IwMwef02X4/HSZN
IP4y0FB+AXIoHWK+C9XkL0+jFrVBVPvTVtmZSpqWwAe2jOpoLGORFLrw+Heim58DVSKeJzdupi8i
M/U6FX+u1ndSyNAun+nQS27n1kgZtDr+s+MlXZMLAebc3UZK/VpusWK1njN+biT76HX+nNLuReNo
q3UeLZbQUzE3U1OfrKZDhP4ifTYuNOJdFSdcVeC9lnz6mqrtCjQZGNtggHhQh3b0WS+KxakcH8GJ
Clash6IH1y+KLLTOqLhEyBwp634a9rJqHznRpblubiGmEHVKpqOMdIZETz8VtDmRTd1nC7NDG6/d
snbNJ7DGEMLS0NoReMRApdMyyINYhTXGDmNBif/miDU6e7IEMlyYixVPoQruPyYq2bcEevrdZiYm
s5E6YI/Y6ZQ+1q0L/zZGETG9miWIDEu9ZIvOMNKAA2BbQpH1Dus5aeCToc9/QlHUaYrdFHRmi3AP
RC5AqgWJhQLgOPC3tlBdknpRIEoMRQ/h2+vfse6MHQkUNd4ue1+c5bURhZJ7B7kkL/2li1QSUGnI
UlZnCj7OUZGu7v5E8UcfcbeBDEcfdAXTtPYZ5EOZcp5IQthuqFEK+11Qoj9RNjkkmZRK6WbFbG4d
45xXMpbTvmt2QMA8+DoiWTOfhaVQdsWSbvY/AplXy/pf3Nh/u9jb4oWkYCB7Ax+h8JQpDOiEJ6AA
phH1bhZGzFDq1v8K1nAaspOfr5YVe7LRxdZTRAg9R/JXvhGbdpDdCENi3sEQ9/V5+Jrw5Cokb8f2
6IIbyaqcgzRY9O6dPDRbduzOW7jTITU35JqfZittG/q2ji5DXHb/Eq/rBhG7dEEOE/XPWNf3iaVB
EMZcFQCQbmXqjW7Q2M071WJ0qa0rQFAzjMkI15SNoALzvW7i2bEAZbj/PqlpodMojyedeiypW7Jn
OnBWs7cu38Bv5QxvG1IjJGf5LaXFS0K8fUwsfN/gUM4zmjkr35F7QPpS6D+rKYGFbQUOYhn2ME0O
t1PyBIBbfz4CDieaFWvm2lMTAmL6CYA/lNoR/bagGjFtw5bAydEl8FOJDtdvnoyxmS/7EQdPyFnh
REL1EhaAW8mOnoUdDpjhiELhbzd2N+aFWqnXi+Gzc0S4Tyb0eJB5E+7ZygRAM3RqWw5A4o8016F6
2oc9W3SAYX8tvo1dLgTsO8/NAAWa7dpBxg5iI2qNBmzgqzh081I7wxjU4UsvGNlt4swk0webRKfq
2BuI7+JJDyS1OYvlI1zj+C0QG+9FOJLVbV8Yvq82p1lsvMOyMdrFiPoxo/p6J6Hp/PONzvNtsGyT
6h1xW2Kaz1c4PgXXww+mSUV80tvLqR02UMogLI2ZZsUH/iX4KierLPFoLBmPGLjI7XRXweXDNQXK
Dz6rGPA303CHUUU3O6NLEULPIthirrv8ZBxQ18927jpXusfEaeKwCI3n+iRmVNDZ3NiVZp7fpdMI
dPDIoLIEvIXe0J/LF5OzexnAcV31zmhotovSaFFIQo9eGLZDTnO3P3bzZyM41ZkhKq1KGkgXas5Z
LEwFAEOS5iRgfQMhNJvfHqnmPxoiiT3avtRLPeuVgoDN3FRA9lk52PsijI/6E4FSeP8Py4c0GoaA
rIfVXhp+FnI0PbuG4XIGKiIfwtvyXZ7NqZTLB8OpBHsiHS56TJZupzIoxOCHQGL61MroB25DPzwa
KGVBk33Tt6Gb1EINjO6UgelqixCcLFkAdzsSGwRocjE9nRno3ZSuk3/6LhgQW62A++IlEtyk0YJs
EV3Cp3D6T50MSCJkSOoz+gxtcUitdZQo3K3DC5wXfBhbKtvbSAgv0TGjVLAgZEvsFyqYm1enFpx1
ZIETRa+tfxLmrQTe5rC4VzA5yi1Ph/U78IJc+bMSa1LuJeupfwaAGC3O1htIAMFFtC4ND93oRTjD
LVTgTYlQ2Xvo5G7ceR6Sy1891ZrTLYdGmsu4+Axsqa/1uqzY1haYPgw5Ac15yqMIlRZPffxGWq7f
XzHY06i5ksQoyePHv428qpOZFOOJZlgmk7ri30Rj78m4vDR7qNU9etAq3jwpnQnTz0k42FyccOwB
L2mDaKmCE5cJeRXJFQvT0k5qCYQdwLGSGgtwo4igfolkcpPAA5nOd2fcBcYG2U49+utP3ZrNyqM9
yOlKUaE28eeDC3s3/28afqtFHE7dS6gD+F90YSJ057sQMChIZYneFgiYhdhU1ExGzdB/kMEQy1lX
/OvHzzrArpFHg2hKLBhtlubwIUX0cnMee9NoQ6ciK1n7LHACdRfw4EiUdEvjIVBjnXcE/eAoPLaX
Z3SGtwTayIZZsboE+fTqlFu+6HH8Obb/FvGP/3Xp15Tg8Y+vs1oQTDYfkUhhXoW3gAtmU7WGx4Hu
W/8kSfeIryV+XxCK9uLGzHGzwhn8l4RWDJ983jJK06EVFWydEddSS+e0D9UWAxzOPEzIn1yz/dBm
09fIGsThhi324NE3btVHwI25xlvn+4XqXcElJunAG5xp1/oZU2v77tTHtfZA/hslMI0freLZstxq
gSGTcbwACsMp5F+SGovMA2W6oInSC303bgpPN0M32fZqqoPQ/1VORFYuh3njIry6AKCL4U3ywJcV
CJqsIWjo5vn3Da2/zxn0KbRySMBk494k66gqk4TUP73Gx/EpzxpXXIc4WibfX7rizUuNW3Kfgpa1
kaCn3o6Hx7KA9ORz2vLX3kUeBIi0jhlReswL1Z2Qu+Mk7qgyyseOArcuk8Ht+2U0rkDi5fXw0OI2
WyEShivbXG7FbO1jSJc0J4/gTfq4NiqRCCE7UZHrYaWQW91/+OstyMCAtt3ONZdZ7p6jgt5qKf+y
XkzGR0bhZOVn7U+zQelhZq45hM2AWH1zqMYQk0XwXWI63nJVzo2epHle90K9AWu6TVhnoBOdzv4f
Ifv6yLrQW6GwJ49ctyAv7qCQhctsbyzBHVmDL336B9OQ2fuyTISlFbKhVOvSXKkq7PAxjGM8acRN
wu/3xOAFWZMb0tukwwotNeY+ty8oacM5LkyggLmxFrwo352zt7PU+HyfmBc7Y81P+c+0Fi74TxOT
fM3LrvSdB3H8DRCKkX/nbo+Jse2XnBGWG7G4HaXID+aUKBD6f7K5gBNZnuEB9WxjeZDrmDp3Rkyv
8IT6tq3VWFIToyegnJhlEj8CDm65JGAdup10EdPZxMs+iFjEgbeqbpr/3Auk00+akA/JKowfUZIe
aEEUvQoaIx/6K2+PzXiidwYXVrCrINFCHZyIXLpRmeMfykn2pXL8LOZOZpP/MFIfIXMxSdzya26U
eosnKSb4say1SrSyoBvvOcuxCwm1s3VAqL2pHSsXch2neGGj9vZzAUpqZa7SuPrihHdhKWr72iOv
ANTjnKSaXdA7ul9KhdldXqhsDxqoCaUOnYalBd0CWWW+lGBnBJp74A9kws2IbaqkUVfvR6AUbRoT
3X3MtYgBC79H2ali9TszDUbiE8+rhpiz69pzqFLOBUp0/xsMdcOeEO8icutJ4IhpktHXrDW7E+MU
6URJW9xSa/7cWQm32PYVaiXVZTwwBzOGrK2rSje70/3FbeDHsbG/JS6uMRonstWUldNyyLMKKiQl
e5lHdJ41i4sHLZf24AGEFg5qxgEWAkKbJR+DgoxMcwIuizI5im5SdCjY/BVdVy2Yk0HnEkJ4nRv/
OuqM2g/FlRRYxKNtB7PsDVrI+S3IoxgfbfLJWE4EBqrpNZ4qwxqw4XYisgdfAbCBS6GV/EFhMZLC
+OzPRHpJM24QkYmtbOofbpaB0gGkaTnQQybu6muL7mBWewknVaC/yqxI31b3LkMz1s0aehtWzw+C
Z/EVBL76i3XrBVzCKzJrrWZLkCV62HPO5giTJPD43W2YkrnZ7ipQ1brUTLK+ecUfCuOU89ud9ZnR
1hRvTM85vHdgVaOSmK2xDeEMl4gsnk9pI/8IUvSbPYTLnJNfQ26LKOsSpZAGYAR4t3jBunwrB4QI
5EFH5Emk1w3bux/B8mqh50wW4Op36s5oShusLgXOAGBvhyoBpDAbpTrAXt36I5+yOgQr2GUNDiYw
5joO65taI4I9quY2tgpv8Y4GnTnzMWdgS2oekRbrFww2ldjAsmSnTqwQwKcBtoFNg3DiCEd/BNTS
FOkxRUiLRCm2c9uqW5xuQ/iULMzocfn05bEwQxcldjE/VqHatoysCKUGQ7laAzZ77uYAdN8fI6DE
s9QL2LWoE9GiPShV3p+DC/Ze4jNqqZF9n402Fp5/TSUaJvpxFW6NDg8+pdcFVDZfnUCIJWL8v1DX
kDLeaACMyWsR42D8tamw5ZiqmRcb5fzIl9tOqEFZHz8Q7vm/3Ftkt9GqVPLTlT0DcupZxqJfEO8t
sU9VDTmaGyXf9WLlMXN5sNon4hiCAYbdiHadijCmjN1N3Bwf7tuPNsuDPZu3ubmGyGu6HF2lHlq9
8HyF1qsoV6KFr+k23qn6Z5O46EAxzevj0qqxtpUWJfFMRQ0xlsI4e+5rBGHUUml/EUJyUzmnTqwE
BuTgU5WvsEqOyE3Lz7iRcQrbXSyju16gR77056vKfb8H5d84mHzUpdmPVt6hhwA9vBnlAGQwkUp4
4SxdUyV47B1hzr88LvcbHvvCNJoSma1HJZ25wgc/dGftqFXZG/ck+iiK11gYQ2aOBUkF8v9Ip15j
XbrNZZyPtEfTRdfOPBQSVspFkrAHdrqtM2dU8S4cx18sp4KDQI2TguCrodXs6uYZ6KZQ8nIoO+qH
dZYkw7dhmKibbkf3MxbDMEs26QipgbtiBV7eDPjkMPRpVA+R6oNMKVAdMii11GFMkd8swDIJHFW5
RJ6CWL8XHRnjoXbljBxnLkeGMKh5mcP93HwcxLFgtq2VxMv+rb4oFoPGvbgAVWM5cXiGKfMXDRZZ
AMtm6JW9jrOR/HV4gbR/vs9d1eS8QZLmsjk0btoineT8nI9eUrnAPH1temLm9X5W3S+jCOp5hUvX
QFvv0gtm5/+nCjTkUuB+d0N5X3EfpoYzbR5+BPFta8Tm2y/SHZvnB4BSszsmir0lK3tU9JjOcSPj
L+pZhL7Mhyi20/WUA0LodsoMr0nx7M0NDZ951txotrCfb6bsXSNIBr9wrJLcZd8RqwkL16bk1v2g
2pWfsARHDEaAZdEgu0nmFbo9y7+EGJoTHato7TTso4EaFxpJxh8eLQP7uK1ZFizxOF68WB8WphPa
A6QjkYFCY+y+QNhTsY5iQ94o4HzC6V7QQg66Y/2Z3Tg/nZlLTbDeCPqx4WAPm/7ETzuEf+IT6eFb
UISODsZM/FwUIP6BBiFBwYp2SzcJdIkt2Gxv+AanInrFl9NS2zCTDLQeoy6usgiqxXKqyYSDRbAE
ELb9aNbeB/5Ns86XFtIWvxcmVlYTGZzkDVdlwa10CA/59YJfjgUaUA4xj9CZiUS+enKQVDy3pnIz
FY77KgYvjTKqCuZaybtt6znzy19DPF7OgLjA8DRGqFULUfR3VgqUlsT7r72O/FxbRuRB9Z4EPAhK
2eI+qKKcs04kZK48xOl0by6tuEvcvW9c6MJV2sppPYycJoIKUc8+gzUdW+lpXnMKqzHuSNCpxm1H
J/pJfffCLFDtn/41LpXxh2ti1sJawkayGrGWGbjYon1vEJgKknINkPDnh+8RX0IXG6OPKGFwaeUA
9kTOmW/rK1N9pVkJK8SXxGkpefoEdId67E64Xk3PLfmyhRGnCYxzetuuCV8ru1dqa7SFBg1b6OEc
9EDEVFU8qk5hWIC4ZZw78tQLl1thl12qXu1Rxx3H2lUFsJB3vBf6v+jeVljkgJCGUZYDZWyXtPRi
dH2hL+jlRG9L5IZwuPYUBCXlUGtK7aquaVAwTIAg+8V82p2wLyXRjEcpsEiHO3L7jozvQZlMOLE4
QgyeqRKVAHzOYPapij/ravIGfCs0/YLRByFftFYd2D2YfXPMHPU1geVoOLjCyhITFDnBfWTlhJ0V
UTsMY871NPF5irC9YRhLv9bkrKQ4NUNwkdpzebAFXedMtzFKVbKs54PNcnljrsiWVybhTvN+d0AX
HrnBs6qDBYr+hx+E5DZ1pz7fqhTJhw6lQ/CxFFAYd6CdLZ275y+ncevqQYWQ69QHkN1Oa5S0nw6C
ifpdPZoRbpNZdFznOB1APT4UhIH/W0XmRTd/+sq/8GmVJ/topHFBg2HnAdNQTxw1aW9cwYTa3BXy
L6yCFVY4R/4JappnSNYP+9IXtu6yJhJGwFJWiqxuHoRMUaZ/+9u0mCwj4KTXns25waN1PJqOrilW
lrw4ZjJUXJI/4bkIvxqQGnTI0mqsyVKF0EGbvOvsXucclpaYviT1RvN38Q3ZO+7/jmS4AXzv6F9I
8y5itLMNndkhTwO5dzPXvYl97bsWAqanldwLxPmPJ+wEFnIMEJQFq8Aoos+rCew1oiwTGveiDMO1
glDZGkV+TPpOF4dfyijxltr4DsAChb1AkdR5zXIDXpkD3eaUfFh8Nta/l2odOLhh2ZRwr9Rjndao
a70rVTvTq/GwYxEiNoaUEe2rEc6s/+bkCmGKGKdSkLDB4lMr+jM9433pIJqeYcQW7XSgB5+he5dL
8lnGXLMFy1umPk6iwC1bAiKF++C2z/bQgbqDY7NPdaz4QziJX4HNQWoxZnfLDmtKz999BlFWiR0T
SAPNBKTO93KMyOAtJyjJmdSWnyW5JhaSRe6rWtk2sVChOiY/LNY2FHxw48krx8mRlxeLpWwiVYsA
8uHddK4xjzYYC5TXLT7rDOp2IuXTx9WNcoGDfRD3emTKxtJGyHDKEZjMT3AnqdRJX/vvqUVAMmhn
xpZoEkTDPDCL1hW2UkxIlRpEvdj1LwQwRKD//qN/W4u0fiAeRLuei9j5VLcv97u45Af17Sdz9Ghe
as8borWRTpzJVT8EX18DWzFX9wZ/G4mwjO9y8cuf5eTMF0N3BowH291y8iqD53cincolcjjIzgPb
o3cifbgFvUWXtEd5Qi9KbgdopJxuozPFaNLMlfqZEjdq7OHPZJ6L9KQEUEOuOncE4HYwwWsoXh2A
uTYk3nXwisS0aiPnBD/pctp8SSqJujA/fPqkPoBeyH2cQTgKVHg875ABfanbS7wM7q2GP43UQE4t
idnKbCeGs1ZHWxLHFI0wulqEQ9vgmuxiRHbdOeuGLJocIWOX+/m21Vu00gl4RtD4DNCz7WENBuVg
WDG8roHUo4OJ0m8s0LXWLdfkqhGjhbQjkz4Sz7LbjFjk6NcrlZlnQb3gFMK9G6dlv0fmIqvY8/ue
3GHHGt5/GZlLjrSwTjcrN68Md4bByM2+ljMgCBi3yFO5EWO+Lhd74arGh33uxwFTbvkBUsbPKmKI
ZBUUR4LdI5sYSPlH2kmoWPxPoE2XinvyTXp61hySu3/iVgX/LihHb42xNkcFc3R0sYqAUAKoEynh
gG00kdHKhhVzWQkite8u27rZH4olpQ5vIBQ4LbdS6YSyg/FtjFnl3WThr/94MJsauNmBXEPCqVqn
xTjU+t5LEMzbfY8Mo0rkQOUuOShUMqinvpqTT1+WgwuI0uDQpzmlSnRdMPN5QUU9+D9SEEYtcwVC
x0IhM4oam2jZg67ctLHRBhH1CfQG1LGRTE7skw5R+1IOYdNpUpJrp3kTp90OGERhvosBxY3C9Vol
V08s+RFYSboV70cMtglybujLeXNx9O4bEse5BvUzrUookpQJs4QKR8UPPO0PZlzbLvpCB1nDfX1d
A4VFKxnwsVy6rE0rHQXVMedKtKzs/9YKBsZWF4Ui27uG9cxxU3MblIdKhSOipdC6WBfoB2MWLoEO
hAH4dmn79XlykAs7czJES1n/UgR8hyYqRvsWEZCL+VNmsO0q6psnKpXLW8arg07EYMwkO8bYVezK
kRlMuSXkyTkwaD75NSQiVUPgsjghnZm8A0fxb8R7w+16zNb2gIm4c8WS8SaZOyjQqM+oERaxDMpr
wXUO9LVxjdnT9S69tA44tPQAnmGdnNWCj1qYHY5S9XCRS+xPtoZwgG0YyPIXMEjJJxVCf2CXDNG9
U3hTKZiOVJvH0wncHZhxord2LIORhmBQvdz2qkyk94yEk/1aJiCfgOSj2308ejhxbt4U8W75PCpg
bs59qDqS05+PaEViLEda0ItH+Iq4IjyPJoqjM7CDATrbansWsRIxrkbuBKRdLcJmbMzlO/A34uyt
W/kWwRE9kYOMvk+G6grrhKxpKb6eqOu69X32k9NmOqb5LCL9iirHSHL7j97BxiHk/qJ6xxcoYdRm
bXl758o7RgKC3fyrJcnz2z3POTl8ZKqONrPdZKtLyr3mrNc/qUvQRiMfv2V9t1lmkgiNHPaU5S3f
TtcmWy5P37yJsOj1J04qwmFYfD0BE3tejBuuq8pyCVh/3h5Ifkb6S/wGK6ChVHkkKdvfA379zTY9
lqRfubHqePCutpFErTUHfDpy4JIjxOAx0KRMjtFjjgrifKsoQPSwdtkrcOHtu+4oT5V2brVKwcaB
KgCHuNllbBDTYUF21VQ5prvPnwvpHmgpBcZfZsFzXPTs45lUXU0TyH0YQiDsexffsMOVAQf4syJT
pzBsTdtBxA3W39KBTjQl3MoCw8YJuEXp3hr5Qjps7a5oBidh8CLudob2kmF0ugutYmWhSxevUFAW
yGqBD2KZua7FJJpkRy8SP9peyhwcO4wET87/shzo5AV6FoQNObSuoTd6bh0g4R8BbhsuutC9Mx7+
VbIZ0f22tBgkA6xyYfm5EnkToao4nghUsCc7iHcLYZps9aLV4YcORr2lIfcENgrWkhrblDh+MItS
1K6BCbEfEAzS2C7T8u6PMyfXgopTTgXPnpR2DnV6fX1Lz+YZ2j8DtFuVOiRpLZLKQE+6rSlSM0f6
W0xSWID0TEpL+poIb3L/AkQNuHMkKAH+L4zqfQUu0XkkYUmiOu8wt71duNpLAQr+aEU6S+99p6Ip
gupa77esUIJZbwL5pUrlLnbjVCcmlDRWxEupo5W9JpPgUBhhLklAMXXxVEiaKPTTiM5v1riMQbDp
59eFCGqimZsvvnccNlbXYhCs6K0Kix5/WN1N2yWiceKBsmyfGohssD/FPVsMYCBco6cyIdh9cS5g
0dasE0TFzksOz1xIJQ8uPrCmk4PtZnjcDvXrHZ/qvYBsu541qhHvm6aD8vtTu/6ZCdxxzb7trJIj
AvxM/Fon/pGnsCxp1jLUDdIMsgjT+mRcbKWCTeFfic3bvbM57oimdxFW0wE6pYIFqSMlMuNZVpPl
plr3jVORikFbq2WTqAYhJ75FkJsfSZbku7phFGr3OhjVPcf6V3VeYhck95ZJW9/x7l/9J+Qp1OKT
lFCvQE3ugT7YPQvj6VNnR4DHqVDDqGvUtFbn6Kqr6I+lDmetJdp6zqG68t9NGT4xL/bFSrrvhJr3
iDnrHqy6ZKx0FVoiT8nrKuaRc+3htAaQPyIy8gfYphS6vxnZd4TTAsnSTTai93eEiB48W/hqxrWL
N+aGxpibBeGKAzdQjpiLClVqTNhOCWmlrGjvE3eus0AeJP9IrbMk+D0xKFM7zPYbgoOpgk7yRRNQ
O/t2ady1Vrt9xo4qucTG4dcRfbdsjTP5b6pM/wpxg/H6lBeC4mSGpFJDwUfsWdVmIocUXC1mCe+P
hAzoBcq6Yu6ij7cuxVZ3/mrZ/JmmNzV88GAfLjQdL6o4EkUFyX+Jpu9kzktd7lgc1SRgoS1X7Li6
o6jeqRRu4fAFaJ867xoFj5q7tCLMxYiJWRbqK3qdKTp5h1MEhPb104fFxKG48MX9W2C+KffyQAQm
PWzNYrlsayLTYWyM1dJKMVgkV0S6Js3FHk3m9NxOsuD5Ek/fK9b9n2AVevBnVIGy3Q0ZCV+EEKDX
e3xa2Ksgd01g3efY3d2Db9dva+Wawfnx5kXmvfx1ij5DD4YPg01rhaqZ+33XrYttIwxgjdL3pls2
vfeUm0WwQIwuxrWHy3qszQQiNOMtDAaLniPRZdAksFL/m7dwXgYzifANiLWvDN6yQw2RWsuKvseA
nWjxcV3L/ihKbq32zji0Ovv9RXYB1g0ASIbgSx242Kvd5X+OvFCJiroW7yeRK92VpmqlqUvENDjO
Z7ic3AFh6YUXbZC8csDq39SsFgnXRsM8ly2cQ4WrYk028r2TSTfY1JjEuoHrS28jbRlV89+NVhHV
/oc23slLU1sx5WkZFpiThxa1FIDqKTImDCoGSncm47GcRxu8TDdYAHXYLgXjPO7KTTVvLj6gj7o9
k1ZpDxunuhh86ZPSmJxYWQ+ITjIIV1QnHyrTp2rofgcum/E1FcVKJPUcItq1eIu2n71V31RVjqQo
OTbzDhKomWKeTbriLECsfIcDF6rWldItTqjgmxcL01HKlOWg2z8vWzQd2nD1ZCfbTXLTDIDyBLfQ
yd5WlhBGXWz5C8z6h4++1vyzKn8T8dINFlRK2qmfvCHzAEiJl0B5BI+uK/0GTPcQ5c3WB/edxL0C
2WRTQZaJJAh8zvnhmVAGwtmY+rWaIQgVHTsc1SvTOcOhV85xbb7svx5GH4W8WCAPXaeVGReNXUI4
2ZruGi3pFsg6plto3wSyU5i+B6gf65SKypFTXPsesihrwbmLr/kSzkRUNEoJHQ/5x59HwB95aNt3
rIcST/WMrqEhb75fWZSyICidMjJhXMSmBeJVBMvZHouH+XZWrSJqV2zb4dGx1Gavas4CFS81XL/Q
7MET7xcrAdjqVxGeX+oFb1MB4fo0Jrfxj27PVFOrc7FoYhIzCAgfgnu8vTWIhWREod4wO8P6zlvH
GUTZ15A/ByAm7bPkqfINrDh1L9Ur++RwhSxfs9Wc5Jz16mqVnimeA69nuCBIL2WqBQ9Wgu3cj1Vy
RN2tASZgqRzjzAKMGvY7YAzdXv8cPgfiegzEYcsmZ+xMu3t8BotPjaiS9BYx3y9z0iY9z9CPYstx
Q4AbuCQezPFEmVQNzUaWjrceOLYjufS7MrciBcF7sVP5X8I+0ZvXRzD0ISX0P+c5kxSflgBV5Q7G
ntSDXfcK6NCJlTFKGYEls5CmF/hp816KFTkOpcYxHaC3BS0m9H4o/XDzemTE/vTCEE9eG+z/9DIF
gTrSTlLdlCqsA7dQBrSyymd1udUt576SCcUoizgNRs4HmvsHlKx+BZ+8TQISGr1v6jXdgtf9EIO6
DMt9kPNN+y3vQjEfrPSYo3B2HE0OGp390fBAy6jSmwGCqv+q9Ml49QM5Iv51kc647fSV4eQzIJHH
//OCJ2mud4o6V/6J368l/3GMSDqB2beKVGj9GTyjN8gFRGeBh9VDSGTlLA/hoF9Y0GaXnkFHXKD/
AoseauTqJryXerxpHI8bnnw0ffQvHjpS2kVX7H/McwOuSSzkvmScsW/t+MgJnx2B+wptFT2oC/gB
baduk+7pEV0uu0JrGhWqE38lL7WL7l6zb6MdH1yKV1He5wwA5Auv5nRyUneuMzihq0YGqSBDgiUs
olrJCE2x3F/eg2iuM8/lmAbaodvyXiM67wGEEDmR+/UiorFOd+UEpT+aKPsqacLjYI5O+p/xYxzk
azKxHdPz9BboEmSskYa0HcJOgRFdHIZlHifMPS9Je60t4shrdYJyuL3Ed9nfvrWEVYPhcp01LdBr
G3064howdSu4wVzpKVN3sDMiIvj8rbFwKoc0144a4t+j1mfWRCfQLIbKEJ3P2ZI/OFj04SIUQ7gz
1E6jzWCnWweQNTK2Bm3v6Kdlrm0+2rFQk6WaTm7xMEMzQovziFEgI2+uPHGame9tUlC4UynfI9oJ
kY7Fmsv4GpDHEukk+W4arZmqkfG70nJMG/tnlgX+zR2qmepfKGCtUbq4wAkF6iqSU5YBpzkvMWMl
Jtuo/VgeC+wDL5UMq7g51O49Hafv3ALG3VmJ3uwMCKrg2RKzHRaXePO8sMY7qLtbyOd1ZCk89A5I
b0mqhztnEg7Y1eoyuIupHDFzE+QZXyRfDtr15ELHfqbdVgwOcN4hLn2bp3oDeoZaGJHeYrYkjmAS
82fHDtEuhhJxZWQNO59Lo3aOvdbgbGkT2KSr2Amty83n/VM8gDLSt2gBiXM6mRQPkbzrV/UUvrrn
7NnsJw61+Tsf+13yC6SpNBpUQLZGDlxprOVhD+e15/klrcL1EmZ/Zypcj83oElBl4VxocwIn3WUo
if/ZuTGDJyctZRZEmtb4ODa0iNVvdTL+yWgQOUoX/mJBvDmuQ6w2hOOomU8cbtAKRNw+R/6XqjJa
43Ct1SGrgf0vq36hBPgKR78r8nU0dZJytasXqUsQfL0w4UPV6fiSBG58dsNpcCa9O3NF01KOWh7C
GL05si5gxuOzSD4Tdg+hA309Hf3CJsVYP6KT2Yd9buxIrug7skN2B6FNrnvXeA6i/aNrhyQSrRsL
ohG4U7PrNYGSYhZqt6kqW0iCylAdHg2xJSFKHId4XPswRJqpXZUrJPV3YBmFGNzYSHgaY5Ie1KAy
prG9+3PzDuDkaqeUFiIVEotGTMEkCOmJ0ZSF8uIPGt/pCtoaKk0trwJ1xNHOd1VcT6kqEtg9+Jse
EYPWoLlOgzbE279AnrlJNkNg2jHMiSTfuQgus8PTNihWCTb+kWfN4RYW4eUcx/uYGC+75wayM6UU
H047LfZSFQYfS28Z7NI1UnkPxOfEdgUXrKxGLOGyZpvMW+VWCkrZEInAsV6meHtL4U+mrBk2PImH
DNXSqE3AgzvPfPS3K4hXYgL5hrDJVvzAdGEe+XO+Jpg60iiAuObZWu2HFCnhkkV+Ub5Nb0gGjimR
LWMOLu46Ed04zai//o2h+eV/mqgD2ac/8vOe4Wv1uG0MdokPnrmOW0fw8KmSxUG7z8ixWTgAGkU5
VQ4p7BXgcPJZc3SwIv2KXQEyaNWN8RFFmtJY0lu+k3AkwCNBxaUfCE//o1DXrNsPU1fkl4Hi3LTt
XxjJsZzl9dogNbYsXY09O/IS0fBiHw49ZD4NnkSeuXhpa1iWTiLG63CKG+yXcz6nb+A/4VwyyzUn
iS+8X08kjFKcY9E1r1q0kFN/+klGGd2Qlf5mNzj1IrN/LpVED22WpHdmGRosErIRNlu8J7renDjK
C80CO3krmBLUbWcf6k32GOyLDdpGVO67QwcW1npNP/zwZRcOD3zGUm9nWoeQaOH9nmgnHSpCnK+D
ctbJDOIAvL134wEReGutWVV55morrJljxfkVFenIiA9hvmZzP/zdue0D6B+l8spZELGGE1bby3q/
SgUSXGU/OBHkdth5OTJ3he5BPStdvEEOA/kdnaKalNM5g3Gux35YvLY3fzXvmm2JdSav/X2BJDHZ
dHVorvS/sBzQXkPCTAU8OHy9y20QQrediNwUECtbaYNGb3oVtM0po0j1XH8G1mlRLFNKJ+x6r3zF
iJ5xLRBzZELAMncwbVmmoHrOmU1lt01fi/0sbOc0SjHuixgWglp2ghEskVB16IIdktpU1PSYRcTH
dWHq/49OAd3HRbl3OBTVGuCJvwJ5c2PdaCcj88Z+9wJR0Al6bJlE2I6aRnsXnLGraLO4CynFDGtM
w/X5ryFbDC+7HFMgTrpbMghS9O6s6XordRgbHl+oNgGhLju0MEilvj3xJ7McwZEIbup8vylLHjc5
JNxlpWyWskXmuEYJlX9X/j5JZUNNoqwxIWYvu85BfNOgxuWgKwfi6WVs1fZTHXrJVVNrtY24Dkp7
4r2GMrjC7X4236m6OzFnVJW5DuXv580CEHmTBOtQc8SRZq0V9PSx/8yUwAgkCy4ePr+6lMsotKab
hoU7JdbHfsjguyZwVP6gguqfISRPMHwnV0byJ6M8n9A84+udf62IqV+WztRg1IN4ZBTa/bloOPhC
wJjw9Na8Kbxp7WfO3pmZPSDCudd4cDqIlDBwCYVvMMu3URSkiAGLq7/nJPNJsE8kGdyLhT0J+vOz
oDUtmyjAZjNzFLHdmgQtgb9JPjcg0tOwZI5Smt0t+Stqle6moI4uAU3eKlS83H3Auvq0ya4TAcc1
Y6r8k7MGwdi67jD7zWMrnk0Z/dFKke4putOoYXYUALOVM0P2oPKCjFXclDcSX+joKguZGlMl78o+
NDwITuqExWLmgMLtSLVXSJYyp8AjGu0AvJZSXx9GFqRHARO+ggjj1WWVVLkqnhQfARbs61Z+aE0W
b3opduODk0HME5CuCFbkgrJijgi3W2xNKontX8D7iIyAG7g1Mpe3zemkQarSR0FWUVFKDrCwLckv
JUzkZNfSgtLzyCQcAT0BeEAnisMKSvVOS6nnf8McmaQ/bIIFKO5St9eCG87ECE2W3wSldE4fPvhG
eDOC7yAI8rNBLS98sWGTPCCS3cOf7vTBbZzjHB6O0csp7M9rmlRNeYWyIXFQsZncdJIsKS+hSU1z
MD/+ymKw7eNHXZLG/PfPXtovYzYZRJn16xxnrswp4jTPH9yhSjYaPjg8znr9JZYKkfqTwqlyVmqi
AegW27AV9C4TdppsJXsapRZ+vMd2eGpQ9CJ1nsGsxDReJJaC4pKsV/hSH9UDw707zQ1oUQuKcjdb
e6JaD2K1UNRu8UoCRXkL84c1T07qTWa5gCVwndxvOnOFswMIdczxPLlhXRc02BrauVgwDoNSkY6B
FFj5e7TspeNYfR3i87t/rBimT8SPRj0TCQipmS++kfliG1EtZfpeOBren/2PHY2xq64nd29nKDZS
L/h1fydfjEur3gLMY+/dXS6CACb+9DuyUDmaCkeiuAso4+UL313Z/xL+wKvBuA71aMNV9Tv+5AyM
aAoN3MbVZq3ZuyTHFKQ0FEKjuHtB51hiGXGeu/Im0+ze3dtN9J7tGBVmvOnPYiSyfYZJk88NgJle
Pn+v/pYnbg1gRdDFhLgFAtwExJzeoWaGwro97bzMwKA1iQSST97zw0pgxPLAhzB2SZ3FMRXPJP97
wvF84QDGE2AQ3tUidTBLkSIcSxUIXVEO9DSL+yaeBZsn+9B+mOIoaTS++wwn9/+c8Uhoe4GYQ9pd
zYKS4FxUfJchwzjOdDlu7KIX/khx2TC+LGn0D4zVOIE45EtvkYN9pvjHEVB2PdnMCdvW6Y9vsu0v
XPsmdzdRQSGORD0vHrOJNid5afAmsupyXtD248mKfFppveHcOF3XQHVeArg3j387eASp+ycrJiuc
IVJLx+Hz/cLIUH7DXlG6SlS92ZeCW/wIcRFucMj+LtvsXCY2ejDtulg3fgvDEidZaQyVkrY0FY0b
/WikVnkHwXN16pzZYrUQ/qkHmSZ42XH0rtKQ8iqSXVTdrjNq/3QNUAEr9ofbDZlDajDNdQn84GzG
cMacIoaEP6tI4Sw1fqtQ2ttWnwsjqmeonCMqRGT849FGFT7/+MS+jqOcohr2N/J/dsujY5QWLLjD
uLda2zVwwU31+WA6RRLnjduE0bOtJJiKheG/eYn0FCcdQZEhhnnMkrF2YZlCwMibVfUZno7zEJ+k
6OYrnAn5BL5Z6wRbOrbomA1vtxAdTm9Vltc/M2tXiBuAdOAA13g95oINBXSXJi8Ho8n1XYDQwlMH
pvIeNouhh+dYl3EX0jveDSSk9sIbz8cSFTuxtyjbMHwuxdBnZUWl9MZnP+N+d7bs74FcE93Y0/Cl
V3SKT0Th37iFFrnylvlrD84QM62xpbpREnPV2D9kNCUj1WXqeiYSD+dah6eJH+Jink9N1FPOCPS7
SQeLnRFKdr+5m/Io9ztVDhngZxtrV1st1ZtxdjrSPSzeRp+ipbq9G7i6OoR0AziOK0a/GwIUM+ZZ
N1b4X6+yOxqz8259lmrhoUjX7jS7OJCU7RiZFRtO8wuoENS0PT5OI1gAoIpoOy37l0124tGlYrzx
jJgHwJGCgon+i0E03ReiIIGjlSC20qjsI+piFHa7Kq5x2rOub+41U7cxLC+bopNEhCHOiCtsJNLf
dmb6bgMpBtB0lC/MMaleLoKb7NeTElMkQT9u7fPGINuhaIhNz6hSL025bMOKdsx2om/bpYXv2QW5
Czq7IO2Vi6GO38lECHJ523vPAqeTXsBHnckW5uTNHYSnsgXj78ysTnu6SRpY80KlAoifWVLtivzT
G/iOuFWzwe/qGZwB+EmG5lIrqtUcXJgIFoNxiNaidMix3iW55aEw9JOAnSXYGrhEUw+M54JL/cDk
u5jcE02BtVXeQ6AnYtdZHVnY65OTv6CLQXCuM6zV7+8709LLHqMgz21hyyHuNCtkXuqCVkVDzh9A
SiB4w8IS9Td9uXdUoo9RZI7I4Pd5T/UdfUNO7jGoUPAt3mS894zSnaAEF3gawr4zEQnzMH13bjWC
uNp3wcJm6H4GazwNmdifiJRrfsAzlAAh9oHjAuijp09NtliWKjwgO3u4C9Qun4zoSJsQ9Wx2oei2
wkyo/dNXpeKYzLMN1H2yByIaCxmhz/n/t6BYGQS3/fPDubMO2LuPpB2cIBr5m0V/0oI60E/wn3O8
cuJQAahvj9cqh/QX4FH52sGKw7SS/SOGZSj8GO1iMT6iFoQWAfxfQLRk/0V1dfpdrDVWXX58Q/uh
VQQL2PEEnd+rZ3VJoHRlfCs83MiKyLkT2DRxyoMXrPRnofr9NJWiG1OZtKqHxFitUvQFN44WogQk
ewsmgMu34HusTfr09aDskmD111lGcWlPQj2cJXN72XFtdt4aXY58WRujr8xrsqBMFPG1up8BMgAs
I8SS8/3Z4zO9TfLTM42MLXCuMnOyLpMfOAQLG/MzfxIXPGLlrh6EXNA5WsH/THD3hUzkKA24dLAI
6B5ZymqL8t6GTm1DC6heHIuifuHHN5nyewI3tAHrcKfKf02avUT4ttfqo65s6AW6AhRWgNbVWdZ8
nuIvkGugQUlpy+azityQcF3XFwKjHuJiijaQn9INjLNnr1bNk6hijfFzs23DsK+g0QAPfl2VzrI9
ekt7bo1TaL+H5keHkKs3gBHPJ2xLtKM9ZyIZC3WQwzuqXclm9FT9sK4HXF+KElykUeztcnFlz7rt
cObidlwurUvecL/lGRwH1Q1jByDB+vRRWQWF/8BRNk1BE+/mQL2BayYgT1oJKDSCZcSPc02tOD2U
QWWB60eGWxwpmCXSTBampOARPK1H+Fsisic5elwWzgtuM16uY3NXw48AwP0lmAJbJX7FNl5LBXY9
fs6B7EgCjYPbXdqw4GXQBSRUXhili9nw0r8QZMgr/zvK2jHndjWSXBkTDP6YfzDkuh7esFHD6JIu
b9oP1I9mKLpbQWv9lTYktoF6xW0IoJfmNkSmFtaOp33JJTIBEjM54iMhChQAcukXo85TQ9fwj3Hm
hQDKjw0OH51hyLflWUwWRi5qE2iX8KJrgdyYMM9Z3+N1BeMQlWS1y/POqSWjs30yRMKmu0yNLgMn
32bYq2g0nNuk4x1PA61/YEYQfGe7BIdtsWG3vKxKB6JpkexcGFyD7eNljC+uJeh4J6U69c9q0QmW
1OaFGj1Ukrkt9W1pMkOt9gxEN8EoMmdgu7I2slFcrXy5tGSU6gmQxYENG6fKeXtTUBiBnN5AApty
9QKa/oDz2SFNy64WuEzo56h2XJfP/q7AZbzkTibUvgr37KA1DuCzQS300Y6Up7VvptnOqLG+QBxy
02pY9OX8q4M8ESlsHOtSgjUrK6r4w4YHScOrWsrm7z2xJxYyBX9RwMuP80PvgH5xTUb+kwfKRgSV
tSoAGnFytRncoW5pf5IXeKEH6EY13ghqg5Ug5YaU/kmSQZudbR9TOYphVGHr0qq2oiyqm68fbg7f
+IxN264y/rNHyvJ0ibERvVTvuLEjdxcQsHDE9bN7sGoPOY9+ml6PDAnrjSV6kf2hKuaILbo4An3F
GXzcDU093J3/K9JEXKLpqhw1G+CXGqNW4n42LuzGxcG/NVn3HNSOWXuWRScZliRSmpxh+Ozh5wQ3
jdgZsmT5Wvx23fWVukQ6fVrHvMBo3cX+FOHs9LzjR4xRXbXYWcPgHTl6SJ7U33WSMiifZJyAHCHq
LQZ2+0C70N5ascRpyEAFY1Cyp+FZpzaKxM01exjmeWZvxgtUG5xfWVYp0aOfJZQRTAXSi4PAi++N
uy5p8WKsslyAo0dTzNjtPCucSfbh3lZ+Dk6/ihB/agJ5845pPygHInzQLBS1os5Jl8ujo4OmXV6a
jw7hwqFl0xg6gyfTEW7ypSfZkm/0ExDhwHemEOsotc0VK7LWqbbIcJ4YhcXqvGkR7CafBemWyt5F
CsVKwfJRarh8YwOQXTPho9aihuUEvBpI0LPI3ePKjUVWoZfsl9+Gxf8OAE/maao+7zAlvUU4jb3Q
//7yX24FPxa95yDBXVgYpWgs4WLL6fVNPG5PZFKixMWd7qkpM4nKK+JxX6SrEytZGN3RQ+N5uP+O
PxcWrWkQWjO33zdZqNldKXdiSpetlxy6RgEkaeZ7pW5ugvA4WIUwFGr5pLBZx5H0Dp4krnQI3oGq
kKOSBj0xdhSM0pNWHZ7ov6TofP5vxR/xBwqAbUNRZb+0a6ue8UM60QhDPu9bU+ViPPEz5LT9+N6a
nQLc5tapNWG1hfVnlLtJx9j92LEkUrcV5ChCd6IcDfGgxUsiuQpQkoQl0gZngUPPTN8Og1UzX6HP
j/U9D+5NEc9q8F3kT3wmtA49saXK3BmtOguVbO/4VdW9wkR0rs5SvKUrZZXPgnQQf74T4JURlfjO
bdwHO0cl9Gn3dCxRO61dRZb20cHcPFGq5znxhJj6nIX6DUPvZfhgMVvEy/kQL3tSIc7t/rteXnz6
7qd6eTm86M74xFzAnfxlolJmMPxXyrRNMAoAPjF8dFmleoGzoT4OtIbDQmI775TwWC/dDzaDDQfC
Z4ej4gs7/UqkDVC/0IBoZxYYFi6FEu4w9ZTzWW48ICR+R64zzA4yQGNQfU2sGRY8ezpNj5Z7s7OT
Scc923GpzY6scV/qnPeeCN3JyHRVu/Muh006nR9uJXfqndZBKA91SAmHJGb41/1XfYGxy3Sdx8aj
yNJRV6+h9FDOts8ZiIIJFSz7x/tVorwxxn9TZZLViNK/qk79XR6bBBpZif+ehSwnU0FIL2fR8jb8
wJ+dHzpdhw4mAbv9KwCTQTxMsUJXooYrJMMmP/iT+4czGP5af97bdXREgAmEyNtjUJiw7JiuVPcf
Ns7n3OqYSk3VQbrqAEBPouc3sMJxUnPSuGVVerrp9LDBk4Q+3Q8f7IGhB9At49NSnm5SCvYRZGUm
0/an3j5pgO8cbgYdPz+RtqzHv3IEAQ25aBs9WqsPAtiUaEvSveshvlScv56tJWqnTdF34amFCsNW
iEAZgfpHQRKRIe+aO/QRrbudlNFJqBZY0o4EX/WNv9IGFy3xzQLTNIshqzwU216W47z514bUApjZ
Jeo8M+0kIU8eOIqDLSCz5meB6fdkIWoRM7Z3XZne2SDLbbkmjiQm3stfWabSpihUAqWQRLBLShik
CtsHbmkFl3HgnUFyzqWzSNp6SkloqrqcYptuXniR4ZLm9N0V024VSJobLZck6Dv77+90p9Xcn6Ek
MMGm/H0iMqo91FodCbSKZSYSUbvMbIEiX52st9fAq7K3oUZWm482JlYZtNkwWD4tZRHiC2z6+q82
GpiIBDX//D71VwfhoGEexh7mU6jkSBcZ/VFxwPtMnRXbComGnqfNDtoyQp5sqGOMU0XXjOgLoVXj
FFSENvfEC48DxaLPAi4V4z0ivW1BGzU8mqn5GCJ+KormFirewiYA1FX9nXsaNEZjCZE/ybeyIRAE
LoS4VE3heXQsVHxYZSGNf3lgWX6C9khBO530v8FG4sNs9mdgZCN/dDK1csYqxD7zzJTb0E5SccJP
AWvPJa89yWJC79ryabvuiF3nMgyhczqwdvxgc2Ga6qAQALsrBB+kjEqSV9giWMWf0ejExdS5r4by
EXxuLCwey374U97vJx4QDVEUJrY4feKZnq8XZMKb1GLKf7YEK+h2XRKQqZgcL9qL7tdou07MFRAA
IfreGcmkjZsCVUoxpqbzC+Us7SjoNQwOmBMnI8Jl94Sa6D5VrzIRq726FvBD22ke0KWO737Yx4U9
pCIZ59CSqzR1zAed7qZgpHrc3qPmr/3yybiIIdNnxjMm636gUaDSqQM4PPq/89TTAA0n9Y/SWN+2
6cwyfJqYnlT+WYjDhb3aLpLYWz9++Fp932RWkd9OBNYuI3mjecMPROz8MlEqp4Y8LGuFw9N5g8vB
p/YzRHec81qHlU4VEXv3Xm+P8q8j9L+fAwMDBQrXpkRC/56iPdhWvt2Mgv2S+B5UcjeZqdIuVEMR
CyMk+7y4Xwr2xNloVlA495+noJ+axyDQoealZ7eNkxUs7zkBuuOnu4Vh1SgoRYjL8h4D9EXZcvF0
krGqls++d3wxrtQ6uD/G4q3FnzcqnjrxPPEtHZiAIxDfdM8BuKNFkNeAZydS0GK6h75aBlXE6sxG
OYX0a2N9Ci4E9nVeJQ6cnbfWh3bzZ3L5vOn2KwWI43mkMAcDvMl46jh61OGtqrpaux81L+XhXuaS
KT3OI67k7Q1FP3HGGJ/TFf2fqKE3mcPV8/e1lIxhCN0ZOld39wB2SMyjtSwgbF8akagi5IMUQrfi
vlrR2BPmS+CCDMNP+yRAMqbnVxj/pIrtNxXJOSm1TGlenEH6dryrEkwyEGqX8OXZuQ7vgHZq4mo7
OpSRswhDdPK3bwoWqQEZUQ6QqNtsWfQKIJlFjRiGnWJKrglSzvWPbA+BUnLt3YtMO2FcZ36034p1
u13+xiJDYZuT2Lc87vUuoXDNWCdK9HNCWyqLmjz/vls+Z3WIHu80Tjg2w6i87KqKS+9dX6tyjErC
eHM/3bm1ncpAH7SOKIRYTbzqJ4tiE+I2lQcXoH/t5qfZkhxpCkSGoekG+ZIgPRWIoSsyc5B0P3nA
X+7vwPNU2UTcoOGWQEOH7t4adyJmrTx4hQHlb2KTFom8XU7dzz5IdEi1UmKBCvbWn3nHfd3d4U28
4S9B4FBZy2KY15rVccPpoEy5NvUrQ1fxQ5s4m9jS2dAN/WAI+cVAKL84Caf6wGO8nrbAQJ2CRL1t
FN8m8eVwN4DzdBGxiaWyRAgt4LNsHPHsEc83tb/SWOTGGNV27/Q9ZJWIyKT8wvflFdMBjrRau4oM
N9VjW+LwFuVIZO5JdzDo1tMWZbqp78gRGXX790KIIQ8QWker9TQ9gh8VGoq+Et3ieTYZE4dn/ssE
ENHckcQYxSbY5qM4DltJHYOOsMcBAKLjNDu8Zc0VnOse48qcrZPTMy+AfzRudUlqN8At2EDi6efE
tmCN2wWSCotylg0xa42YtTH5/Qx6d8FMG4HDCLGcWl2/PXkKL5VvH7xPTLhE9Ney3qF/+lhHIt7f
mRHtLhBoEdvHMlIEqD53/NwUKuMV08t52hWVfjqOgHDxm4XisXoJiSeIFdC2b0VNVpZGuAcjbNyF
MeXSbZpBJ4EnrilPgqeNIHvv3WzdVO5f2BRRdR5i+s2UXYPz/iAIKnvE0Ivevnr67dVGvmqWU+SA
oyQW8mDzDgnRbSpJUdsqNEbVIlXgcCqbCs6GBGBbS3NDqbX+BK499bZoQ5ZwPqd6ch18h4OgN6T9
JdQnjTg+A7DykZMeQ+W2KRAJ8RSy0viy8ji4GBlySGMWhdbBqSAFsAhWMJhucxgvAHvgjy/Gc2lB
1jQGNPUA35wz5HvtBRZsgPnvJmI0+KVv9qNzPhIq9Jb40xH7U4mPneZ0p/Yvt2Bau8DOELQTuiOd
wUi/Qb7vhwCRZOe8RrpPob82lW18LBlbDCuI+t7+uvxV7XrEFtxNqEDtHVxq4U3nyqupYp7ngldy
Zkx+pjsPxYja8urqOlGvYiOHCdxNzg3kveCHdu+HL4WPEKw1KtlV0jMjnW9POL/SRGQoPTOGwjQ8
H1tJu/1Rstl0kAOrbcX8G63zhdX9BnuvgUUzalIo0Wqi/kuoYvrv0DWcz/jQ5mJvzVrI9u/7xnbD
SsvRrCTTZLA3+uWixTNDmRQ2aCbgDDlMA7hJ/Wg7k7PfHHWaebI3Y0w2QDEeDoa7bnupOcii8Kq5
Z27fcbnqg6eMVB+r2P2yac2ykZXQinmn71IvGfxInY8ds6GWcSTTs6xdOLME8YQhqVxWOHSRSMVs
WDS+qiPdWQlnoRd3sAbzvdgKB68zE+YKNNptnLVBVDSACPbUuItZWkIxTuGxVvIuk3JH0DYm7+6H
H07hzqeVcB1y0Fzu2jnU2ScRU+ziVJoqk0ShDGbMsnWWtXTQu8hskR+b5FdZYBLf8l/832ctM7wU
jYec57aijG5uksx8y5uTZifb294RiLdxGQz/yP80V0xgawBOi0isHELP1Kb1VxAXsRJl603D2nl2
BcNuHrfApZs6a9Lb8BEqz7ft9RSvWSMEodKbNXiNGXnaf0U4jRwbrZsMEceFG/sfc6ck9qz9QSgp
itUB/3M79zBCT1q5zf65COOyzum+C1s9uqSHRcNG7ISZkZbLy8acoLlbzCCVDaOWLYJbKc85+pAA
zFeS6XawR733lbPmGO3nyWDDThhqghz5RaNekYW7/edwEKIZaAuczOVklyBzohK4gcfuFHPlro0Z
j6AN1EUYMsC5vmqtf0k5BQ8uXaukbjL7c6qqQRTUmknyBqVUmeKDghxfli7Rc2quVmUHQ/gj/Bg3
tVsnUZhdAR4gaJ1tZK5sMX4IyHwKULq4SWGe5o3NUSHt40rKglrB6Dj1A+LrTgps0JeunPJQzRgO
3ZeLNuY8oRA81mWKWOvB6nbvtRYuGArjW2eQrTL7C4UeHuTO6CK7YRoJIY3uR0cEbZKMt7br6PW2
GineFuWN5MlvOrunIfe/Czxhh2UI6sidO2SCB4Lb289+qYGUmQtH3y1Jh/zqohaM96D5KWqZB4zu
dUaCkHae6e1uGqa5FDo4gO5Q2gkETukF919UR5/CUrNxDhdAr3wFZi6I65Abb9opy9EYnspHuNeO
ijXFA6XqEJeYVHof/r6pK/2P2ZKZ8+SgXB+kfFSEHPwqqmaTOUnUBn769c3LJ4YfLorNt1jSHqQm
4+iQF29H0E7mOXaRgVHQO7ehH2x5coBFOuD3P8hggmp+QcUE8i1AqZc+Qb0Qxhn9KLQ9tK/ZrRGs
rJ3ZxFiDbrpPeKfJ3X5SY4Qk3sUQzP6bBRSBpcA9MLjJUx4ApFxsCGTgjDnXurPAvuA38B7RMqi5
6yT/JkVUWL/orFzq0xlkWj+2l9mGqcqtxXQUTjOmcIK5rdVRkvXdxSZnTksawkxvM8FgLicmq9aN
7OmJ4ra2O6Y+1KaBTCdRltv6LbLvoLTPnbjXsWyaIyOvzI1L81hF37/C1e2rDBlqWXAwaD9zpmTA
k7NVam6QubgF2uynyZpi/2bhpwLQE2sNoTbOKyuYoxawbZC8/OpcTx6Xf1TY24L+dYanaFAmjqor
hyC6e+L79+LhdNjnTbQuVmQKnorgVpX9E2+NNcnUHgVYUHauHLxqsSrvW3RUTFvM9GAuKZf0Fah5
cVd+Yohld4QIIO5h07Yoff3uTJs8ERlLmx44+46uuc3MFnQk5R5RvIAs0oqNFLjdgvEUK/uD+EsY
Z0vb5/iMd8UqN8SgcibX8fOjZQs57+I/mSWWb8mgwfk1DP8LZiVCPGC33bRgA65E/jOjt7O8qGat
InSDM7Afhq2KzhXDOLklehozKqOORQMAYMBUMGkMMTHNoYGYgwedUAYU8J86YDu3XZgFr9RkA8Yt
1pQjlbOjNrEzqGjg1/5vd8pw9t9e4wwYSr30ngb5MWLxgfrUEWOFcIGTpCBI3T59P9iWkOnJR9ww
xgl2QrqaRCpTktbVoNG62P3If2aPpt4aGyhOP5a0wFmJH/DsbPVQ89jdDkwnMwuXgt5ejk9dRYBF
hD+7AkS5JvmyGEkaaYoYIY+rujR3tU63kYNfH0pbVdz+LI6S6/Xt19uaSIrZw7OX2NmZXOtyQ5JR
ANFXZYLwIpG/YbMKtJoVgdJaXN/Cfdd1BuzeW4R7/u1pznhh51G7/lpvOOLzMdGsGefsWY8JumNj
ThKvs858LAL5n93YxjHsgiJbMnj6le3bzFZ6kD6vFhXSDjmrQ02v3HK0gWVBXyD2IIpjnEP2inZ4
aYz1RsHn6ZISTpBzC8fd3ru18OadVYRJHTz5GRMfOIqie9ORQSqwLptMBsxV1HXMmha/TurOZUdC
u3gHtWUvo7BYaZP9i6SN8sk+Sg2ikh/GvB6igCMhOTJvMMx30QapAGI98jpM0X+E6/E8y9eQZg3B
d9qtIE4ujqXMWG0VNut/Ve09KpTB7qM0zwual5EGX5UW5NVZUfyZLsc44Zi1vJCpfSCJG54QY5IS
gJAd665RCxLjcfXFWhR+3CVKRtMQ5vzW7vfx0Z+NrMUXHtI/Xtzsi78KLApBbBzgUhx6KP5iy/YU
Y0m50U0v0fQwhNLwNlgGzRGOFAhYLQFqG2WfSAcvsdQFixlPQ/HjFuC42v+vHuVSndf6YZBCyKdv
yGND76GhXYKkMRRYZNPZ4uWOLRhqPelKxw4Ful4a1Jz1sQ0pq329yfzvqWC7i2EJimsS01zQUsd/
68C9TlXqbOvVgnFlsvoriWLcWT1xDG9wkgTHZQU09XD3qLLxiIEtww2bFNX/Abkj68C4nWzwjJqW
bAugf7FtMhdruZdNuxhdT/1NtQZ0GjkYmwQe6rZxUJnt6xlPagEo9Z2PQPXmLsjf3Mw8llf8GznE
CogJx2rqsdkQgF8hUOVvkeq6wyiLqGIvEqOn1sIgLPtg9jM/2UmB29MM+2J/tp1MaQJd1/yp09fL
kk9F9+ZJWi5oKgvMcrp11j4IkinNVGJWJoYmoFdtUF8p5WqLjd7JHq4n1ysKj/56NJVvb9S0oTVz
wAjendnTkMKlCJ3snmb+qAG7cEHvob4JKBcoZRisQUxWQ0kYLX+e/a+KtAJKw15OP6DJcGVWukQq
nKNqgmhFo5BDSa2sGxa3595y2WTYdBDIXRtHCiZxXOYOXuMP+Rz3UnrYRaIwKoNmWREgWY4CDigM
b5I1FrWWfuPUjvJb9Mglwjx3XejhwVKQ1Hssa1LFSNKPYLVWHt2nJpIkIZTo+u3I3y/4gAswqoEH
TknmlR0JE640+rcmjUosRkYbxhnEwH43b9pM3Vc83b5LEQhr8XaZTgofDRDUeWTrkV7Cj061sI1/
hcArqJUL4h1TZTqr6pfIB7vb7poWgou6FwFLPtMdj/nHRJqa886W6eVEUb+/UecIp9b/JFsxY2Dp
B6OAuEJk2/fhCboyTCBf9yy9gmtnirL5yFDyvgpxeApWUK3JiONKN1Qv7Z+L9WTtOgsyahig6WcU
+Hl7zG5IQia3OUkO1xO05XvH0g80ayw63d2v4eCpHzGL1nysEce43q21xjx0V5qmY74Aj1h/NRoc
aCYce/zUs/v0+QuF8mHNkv8Z/lH+4Hc91ps4vx9lRAozrOasgiXgOwSdtPAY3bb1KfUG/tsIlMTF
0ukABtE0N+LePp/27sH3kamaDLqZ6X4LnNT/gTL16HyG4If0wP0EYaib7r/CZ8VHhGVxZ+oQQb7b
SCHTNhd+pnB4AevRpufqoIFDgsFPZ9/n9ztNFP0yS5TTjHv2FH9RZVhMPR04iVbGUMOb07nnCHIs
Wz+DY6iBo+b6xm/4+O8x6INUQUyKNFkBaOJci1VhMAYxwSHfky/rlJCu6sCmIVhYxkKSCut54k2C
zk3JlMKEHDOQCa01p1eCfzwTpeGBI52iDF1fAMwhNqNXiJCoN/LZRJM/ahs/CzMlTU4wTVpIMyho
nu7Dvc4vI3bsLuEo26Qq6YSVNsjepdSqWFExwb6nJhByO0cI3+LAAx+qZdE4PYoG9XbZ1leRmlOp
Z8LalgR8atNRkDBPWWlLa2Xq4nSxy4gO6jyuw9IX1AqdSqlEyOWyElGjGKA8RfSJATPHMFoQ1gTT
T2Fl6dpVyV0drymxi/3+KWt7NItDQX8eGhoUDIURJX5VgWDeyNjWMoRIGGvO1fXvtt9ZSdnWZjIp
bb0KnzGRO4QLBjnqQPcuu3tX6TrHFtURYzDZpq8uzfPjcX1J7EclQKLJeR47JJs6Z0I1nXzpFI/g
zHCsFnCoIqLDraFDDlgyuZpyuIDy+X/BYamEuMw7+kj9kPHOIvDLBIvPIr3FvPKQWUVgpOqrCaiy
MYh+pHsznhpElPLigZIxceFk1TLXrivpdP8QyUVS8d4oocpEFqsPoroICspf2sRr67160DlFQ0tD
Ekc1kUmJ1gkXcpwDfRg8FrbFmRggX5JGoXEPxadgQFECifW3dSm3yRLnuoVIhyglJnGipcpkajgs
yUiFF0aWRvsqFtskjLWG4cCj7gxmogOPlbTXSAzUHc+X5Jcidp8kMEBW+Ztm/Ck8U7T1z763QON5
MloSd6+I4/1uYSQivx3XjGrIZM/4QXH/NXqgCGpU4LsS0fDSqAMFSZrpsdDOiiOpnVCUaYiSwQZm
1KKF93YnfCOqATs42+F+OtkF9CYcRtu9e9+JcSRt32499Hd+zhohHkfNWP3n9z9ntoPTbCsiX1JJ
nQwhJhbryZFei/MYwFoHsZlkLSyoItPSm7WfMmpOCZjqvQSE00dwGqHhSuJ9NMgoPm3l1yBHEjiK
OeKMLgzxZXc/TbznoVwfIKMAp6s7nC9gA6wFNwipZOzTrdx00Cyd/zTXx+HH3rPPbRdJHUXxVA2Q
FJGtZ1GkKZXOLc5wWN1Fwizoe3AHZAFowE+CTotNOKf/V4dyOVMG9u4lmLAx1lZ02/sPeczaDrzu
aLVxwiayLzIExxCFIwNCkA0wzWYISSpvav9csgvsYV9FTAU5dbRrfn+nIuxiys0bClQRPm+Qesvg
hQwSSczoPVezSQYJmMCLFisWmMMQ/Z39RP9FKNzh+CtS1NhiD5TcJbAecc2rlA3ZqYqfpitS7ODE
toX2JADg3lKN2QektEci17CNnExvGcG5f2QkKW3JIG47Xnz3lVezHgJmc5NMwVFiBAd+Ga3OQtv1
TeQkLXTvTZDOKl5Tvl8OKsVkCmk9/49Cl6IyF2XpQ4Rt2Y4MyCwVhBFpfxdpI3FwxVHVegpQxEfI
wq0C45rmCC7jptQkIMSS/vdsVWQfybf1J+8d/9fuVlhb9c3+tuI9rw9lOM3g6195s4NLHVdxVakT
F7sPNV7iuuq8eO7Ol8eKKf298O1jLJ8X7qwD3me1Td1la6GH8OILFMqwBVoJw/9F7LkSXnz3PORd
SDaP5Gzq9txj4bDMhzwGP/8KGtLoMDYnd2LmuLiUIF8WXwiS8fx42yJgrhzKr2m1I/prdnlZW68U
sHtR63oXjMuzNo4pUpqh6EmqpwxmB0rgLiwnXrOYm9yQAFNNNTDLZ66KPdOtrpLbGpn3uziazA/L
885eGnLYM6eTNtgxktLLkyPJPC4mWqY6FQx2WCay9nLC+qjGvmNHKuahHBZ5uGseOVii7y1i/F+M
MlE9ax7gtaTy5LvaOjiyxjaWDQU4sTeLZ0l+BT2pQXQZKEKy2+h5ZqA01PdJkcyfIDBfchFRYVK8
izkweDI5cS/tTsj/zni2wilWOoF42vnkt0+kh7L5yKu4wG12XbIs4BsQBRNF2nn4RMnf8un2tI3d
U1XiPA7z0dM7V6Mcpgt16Bc6C3nCwJzCPCPWGCsELwUknIM/jPMtMq3Ads8DzlLEPUHfSycebBVA
8Tn8a9TcYESF0wjp0KDJQeIDCTNmVZpb7WqvLRsJNZdyp9JI3Kfl1rrkUgIRbcGTsd9TRUTfouBP
d0yoaOJ72Cy74jEubjGh/g1+owU/PYiSFqrVpgy/iR/75RflFU0unsEsthilkOYOr7LJhYVdd0qa
C/sVOMGcPVw+tzhnV2LSolswneO7JCqYfHEqS1GBZhQfsYe+ajfCim/yF+UZQURC8T6dgWElqIgp
2ic4wgmsyhg+0MdX+S7o0rkIij2FVJ4nyqzQlIYqbZiSVHGy9hVXEekMn3c4wwYB3XPoUptA0UbI
aC9dnRrThm1XZE2dYcTu3Kbke2LMtzsoaojg6xnXvN99wCVqsDix2XwAHZzmZ0H0U1XE0OU962IK
wecITHpsPMSHE3kTQlnJ00sGXFkksD72HogQpt0cSD3E3sgg7KNi3Dk3DWNjFeUegmPx/30iPL3Q
W3dw1DzllD1mwwC8Qz+sBG3hHSkMPDHJW3NZ/PJIX3eZdgNISDNoPqN0bIsCMwa67ZLEi3sWUTX1
gOnwuSUnWYm+CMgwnNFNAWTU+/55DvmB/i4mPROPR4KrsESzsl5hb0sdeSQDuCt877r6FgCDIJYi
K18rHa7f6YGhJkDYhejIXvozsndqRca4BPtWbVa13m7eVxEEAIm49a/tO1M/RcgST8NgbwTXP/A4
xBRGRtIXMLqN5MKtoMYKxLjf8O/rW+7ebkfkZtbO5l5+5XXNgIfO7tzXzkMIkeLrt3/wez+vJ6jl
ltWZAcrJXShBoVmFCjDKZLnuC29s9LE8RYkOirBdA6rqrZWCcZgoAea3XwMXMQueSXKKP+UwT/94
hEWxswZpNmHxMK/YdGYS3Y+MEExPPPhhCe/LA7hYS79/1mRLHUF8ae8LgBS+5UBH6sSYQt5BRsMv
nFWh5M2ZasWEeF81Qf+T3gp5kNqU1IUxpKmjga//LlI7sKqhlDy9xfTgD5Frxd2G9yKinqc61yCt
7lznkxDMECTgY+mQEbZdWZb4IpdEk6Ud2/Ek4OsjfnuyiS7Er1sWPr2TJfeT0sBoGNI0xyH6dQqq
TWpEZKWovz4wxREXcdnOqJZrO8uM+xkDYlCMFpPsebIcDeaT4tLtiH4Fu1/j05+kvPUyz4QC6NU4
Sa+TdGOQBP8gW4T2RgXPRuHrGA2TVPK98mrqipVJxZYoVxmYfYCE6Ch/aJsjCSiNo1zJCCJZ5ZNG
infu5WZ1kXphKdNGHAqC9t2R9a4WVdIb/6HHB8lySoKSlf0akY+OuPuQx1FPWi/js9u2lJhp7Gcm
98WKk2x6numpxOr/VfbmdH7gPhmBSYQYWxum4qIU8OHsM2PcVXNZk5wroMp1pjOVxVpPra2bR1pt
0vD+/2adaxjz3nUGs62FYGbfbpzy+yL13g8AfYQe0ls0l3iAEb78/gQxoeSXcnq9tXlZtG+BPqHu
n/6Bo0NWAVtlhnRw2a14Fot7wK39y0crws2H+Rp0Ej3B16yFe3iohE8MpCd8pry7e2zbEixgoNIf
Yk1yNIWVKr4hmWu5cg7OSOgknYnt2Gx3QP3Lcd1JhxmetamhzRyFifJ8mfXKPqVjk9rbpsFr7MXs
Enj9hSTxqO3P0aNof0MSHzgowS/v/tTy7Ew8c2nwXOaNZrd72S/9BLYPmfhJDgkfOQXOlPf6iKwD
vn01pgGhY6DGbpSSk8Umdo6KnPV0zMTntE97fMiPEQXOE1xlz2cYBDKQtY3UTD4+WBHcTePU9c5Q
iXKyXFQjplvJEsChTeaZN5IQ7M19Gd3Zk/n6/9tFQDaAfHOJ0kUAB0GURwk7i1BEcbH/qXfE+/iw
/pbwNhLMo1hfcfdmVovI05e6n3fxg9gONsb3equtgr2GHXlONtUq5dYfBIqufV7HkRHb+d7o+guN
3/wAqNg8gzxS7Jm8Jqamhoxp7spD5IJ1dLWLTLUKwsDwkn2YnysEWlr55UuuyZTV8qi982xA93r5
JF/EBdlgLv1z1eFJ3pU3ANqRPnhp33I+EX5SJ2W3B9FqbFzGGctZkV00UEwcZ86bah5MKub5LVp2
pPAbwoN/1nfFFZW+Rs7sovj6eVT+axlG+5Jr4lSLewfvlKvOeYXDOrIi902cFlv2rN5zhDDgfFa1
ErP/y0jlJt47K5p/2pmtlPA5BK5xMlVcyUoAKgmh7c1P9P6j/M7ep0cVdiTxQmFap5xgnEohdQOr
SyF+wTfI+8XRsadu1rHloAo629xBvrvURfUrHaHS/fV2CBnNQHpS2HmQFNjPRFo3bSEHjhe/BjW4
ZEy9LoFzfNfurrdpUNBMCzfZ8x0jz3GlOE/GQkoCGeEiqjea/0f86EFmhMpLJoEC/2aMmRlP0KVS
iZAc/lXsa1d7UKQMc0LJxexjgpoC30TnfocntHBRULcfWrtGYOxA4wweH18QinOzRUAYqETKMZ4v
Mv1BEFPg603+V0kTQArHy/W4fQSFInfWNI+T33EqOTZBHUU9eget6koNfzDvprIXiY+iVnJxrItF
xf5VIrMP9FdRwVSXdEn3T5TzpeGCj0ESSe3ppmCpsZrSbE97GK+vn5YjAbynsfDPlINoLqOhIDit
q5xmU4k0jvEuBYes067Txs3vnYLR3YFkPflnpgbLwyE1rK/Kgtmmk+3ryopiEoZli8Fv9hNG5+cZ
2usG58kPg1atsstPKdmYdKJ2zpbYqJtV3Ij7SoCCEtk9c5smO0g+Y/IGpOktamr4XiF9Rw3UU2l9
bD/r/zQG6Yb1g2vlxBXRpcgrTtSmrGjDadMdN/j2cYaW7X3c/9imgjg6mLkQxlS0AEDl1DIFAasG
U9V/6/dtQyfvyN1a1dmsvdADofk+j804/gz9fsfylfvgm2ogDQ4soaCipBXQGwUwsZj0ZujijVSX
uMkh2mZgTTQFRNPrOkp00MSUrFWGUMEe6LbSRhDph83kVwGmAeJ8owuMc7qd5aN+J6sFKNhP9uhR
cakkfZlGr94RFVG78sksyiBfQsmCUNlbxsHlU0afUGtUHTTji9fVM2dZu/BcAo4CRFhfwxkQ4y0H
RaCO64JKa6l8q5mT5p8gc7VuXFE6JsV9oza2rdm0e8ZuUcFauVOBhN5BGll7tdWKHTm0Yz1qyZja
zDCXUTnimQ5zHA35Ho7CZ8kbTtrSSCXwgyEFuMwLit7IGz+vkIMsFakzSq6ud1VcfMbrlpwMI9m6
83wdTPTeJ0sq3xdfeActYWfJbqCoE4ZSQq86NDmZeS1lexVGlRrpK1nJMNKPX9E9jwhX66xX2GEW
AprKMYl5Xfrzg6ZWxcaEztXaPjKwymJ2y9xAyNDsMtX1OxNPpTLNLOimABQc1X8gJZYKAsEHxcA3
C0CdnK/mdk449bn7tYR+cpuGXIk6Tsv2GiKSsQh/RcddyGVbuGEndziK2i5iUZ670Wf6vfWf5Jm9
HQKpTL6bd/4/DJHobpKBqjRh3RaUbO8OmP04IDYbWPYHuHxS8Cu2KzF+rbeTBMG2VnaouCk/N+O0
8EoNHYVf75HUxEw7Ye2RJvV2f+83TFpMEvaKSOsIZxqITvassaT5bjZFyk9u6MqYVIu7K/xB6t5o
4tdKfcbL/b5sYmwORWke8xwZg+gx147UsKQ5NT5fp+kRdZjNVmwy/z8mGyx52Eg2+mIqhBLT+WmU
Q2pgl9N+LZX81BvVZQXTdi6gLs4owtzSa+By1Ye2gVoJkhvy7BNry/peSvy6wga8aeomt79lfu3k
5UtkbnTcy5uzNS97JI9E8M7NEYDHbYrf55y9mM2zW8XV3MELnfL1+5gSztyiXfdLuM1Ftvsq7tr4
qPEMIFcC6Y3Msi6a9s26R2J/jc9egqbx8oZtg+sdT2R0roHErv+gz7AcJikykJEv7b1m5Q7g0OJd
ofjQbcsQ7aUsw5BkOKDviWFNWbZLn5lWqUepRi+uKIBqAgeCLajPNuMm1qjY+/yCur0w47PBELbt
hyPELMq0sczBizIXOi8fnZwMEbXBmOEUM/ypNgJI5CSGWbc71VY2LxUA5dhuIcxVq8TfDczUX7T8
tmKz/h5dnp33Q2342cmcebFYZ4aaUQ5PTtk6m8Ty3IfmnOo49qsU1GMMZ77EreCXdm8EK1s/8mKu
ZTFOEEyguWlcMVy5oeygFOLiISxE90sYnur0PKFcCvyWWShUMvh3zwnV+yc/Zz0fxeXk6HPVbwyb
IIqdmpiIw0lg8Z0OUF2YqE1lFe+sZ0ydDSQqEZK+wop5aRyNLq0siwWuKKgqjsyGEWMPSO2V6npb
LwUeXpc8GIurDTnHZDU6UPwaJvJz22TTvpvlfZXxOk8BJzlME4VUyYf4bPsW4TesrVc0K5rI2AAI
VUDxl+w5aO7MAspNdUlUxy+8Yho3vbhq8LQhLMBwHrl6+KJT66h2tERJ9AVZzOluXWZsBkQDbPiO
nFrFl7t4Dpcor6+taZ1S17A6ivOflk34oiEFG5WBhYuiZtIoWQb1NfRc5JVx3Ox3brhkJ7JHEKMG
Jmytj4FyU14HeWZuu12W18Uzpz7i7B99ei0fPhDRD9f/3GVYDAjVFahwAtghyawo2w4sJIxutyCZ
ckZvqmATBXxE7Ug2PwPPaLTOP+1kY9Oo5xJY83GiDYU1+zlcElMNcjkdWoCLWSX5U+q4LDbqL1U2
vB11tE5som6AS3aHltHwhmNZbndSJiLpBfWzqn7ylCnX1dnYDus1m/wo0SZJ4dD6ddaBZpFb+Lwf
qpHSfDfFKi9DU8mC7csyNAYjLKJY24qdbi8bNxS9hlpQ0RYVDC1GYN5TxQN1t6Bf+Fp6iO2jBrLr
S+P8ahkP9s/AlZ/iu2OgjHrqxepHRw3tcK12t1vXdO8LHuihP0EqUalOONX+LtPBhSsufIZykygx
TWJpzgYeWQ8pmI6nmLuKwH/WJboQa0d3aQdZ8PrlohdLKf8HiCC4qPmmqFai3mDboFtYX4IF57Th
AAOq49iGJnpPD2o2/iU+8NoO3iiopoMZLQawmkgX2M1xZFkADWawR1AkkCvs6G0GJ7sNoDcPHj8f
9m2yderg2IzbN3IUGgRgUCng2TTOutJ/r6QzHP19N1t/W53XgSympidJDrPMP+pZ+vdye+L78Z8f
DyGyazmEhHRqQR1wL6I6AnRx47u8HNYJNzUKtdI4e87j4RnviRJpK2mlqM9SC1x7v30BHOJ19GAS
cjOcfuVM28mCf1Ii367E5cmMiyQNtFWKq5m26mQSluhmaUNJaW7S58AGm1o7VfGHQXA2NOTaVqw7
Or5u94Sy0r7Ib9p+EMylkQXHyhJBhrET9lya8Krg2AutJzliP+YuZH7PtDJ729RRrmWMiQ0PIw4o
UDJbnbG0b6PwEH1o78pqXlmFW18Tz8QGilMso1nW9J0P8s6B6A65n0L3tT6HFcCU6k4sXTQDNyeJ
VfFIjjz8Hovw5TTZbDUQZrFYCNqK7xC/rN24ZkamET3XpwHvonrsUhvb+0B/0fi0V78J+7I2Muoe
NhWWREhFvAB33s4E2Jj68+eDcuh9L+G8mRbQDrmqyENtLeDom+g+mer++ZM5WPS5g2P3b6ApX4Ze
v/uk7am85jIsb5znNOLnAhm/3tXZAoEvqesmKx4to8tGGSX8EkgXvHiXtIWue9ortKsRYbElLJ0n
vznbbUkXFJBFidE2ixSDz/5axozdIeMzNWkUZczhDA5r+KANJaLQM8fJ0CR/9+laQIsqak6hrVJx
ddRRCxUIHcyoM4vopZpeH2hIMKr9MRtqCPZiTS+iPFyw63gQ5y/FT0MxmY1RIpglze2dX9UIvcU1
HVqs+kRVeQlwy9VZGjcvozqB/9DnWKv7r/WscsYXTDOXyGH2e9v15BG64gvMwoBlBq4NlshgjMgq
2LH9A56yQGZR+bqOFJF8+fR4Hm48JsOnotT5KTSfZeRmLTpXhb1SNKRiRVcK8W2vTuZF0Pgv0G5e
ycdqfKOmjvxocUAx59AezFqI3wg+dCFW9ZC70Zc8w8kdknAtlx1FUjEOQuuwuh+7oUCJP1VZn8Yf
pLgk3Tf7Qf5MuheNRj8CEX7ymHSrIV+ghLNFYQPatYEDEgpKfhBXtnvP4OSUtfS6VxLIM6Fogmhf
LIB268dPPVXEPI6+NdEKLFRfsvacFuk2Z2NQ7aFdGyNfpzuQtWVcddDGlU4c6K4xlgaZrcnLbsKo
0SSGj3A2J9rmzmg1EaPgThuKkE2g+CU5b6Y3vmnHBMN7rRDk5tOuGERciLkYAy/zIujTpFS8IP+u
nT0oSrVzYEJga3Vo6oXJBO+LTyAXfP6Tectn22Sl6l5fivRjNiLEv0l/MkBhNpU1Q2XMeD9+iE0C
aFdYSkhRkV/vZ9gFeNbizx6jQ/b8f16Hoy+END3ZtQlZodzMYx2mVIzPN26g9iwJz7dbB2lfn99K
kRB2sSagHw5JySkbD/rpazwsg+ve5lyj5Hby8OubaTsRWjB6ojI20AFXmZA4uIpFSBNwp2O1RPit
Nr+JjkrfBSZagfkjkjLYXYoit1PozCj8BeBD1GFLEgA3de1PENMLqQr1p8vFTziNn8xIJlC6ZI8h
zPSwSR5jnjEGHaBiE5SSin9cYGfB1rRKnVTpxJqBRk8THBUnTTOjSq5Zf0dXZ/TKbM5iBKG+SHij
6guRTYXHGMfKugwl1xblG5qaDsLfAscdCfKGVb29wrYYF3Al5rguev86bsEaDnk/yPsknWbLeiP/
DoUkCsK2JhKBdQ5si/jOrNwILIOQ7N70CJXvHN2GVux5IeqSL79aRserC/vGndTqFAE8O18C6GFx
g0WuO3zT1isutZkkliZaXI8T5DDr0YFj18STd3ioVuln/2T8XZAuHVSBKQlH+0yBRBm25uz1Jo8k
kS0MfiqVrE4ku4X8ywPKmSR7i0DpwAMpUvZfPCZIYAHoeXwleWFLr10Z4SE1zeOZKIWnj5rJAVcI
XvHP31g/CjxrWeRfACiWmeuNFMGJvDI2EMEgoAhibnGwRhvjuYiVgGy3mZ/D7qh8Br8H2WYPRJIx
5XCSAihwDHyN6MRLqW6jasA8bQYjPHJSCZiS8ZoMw3Hu83SRVJFLClqYqw+8Bkj4LvyrXz/1iEs0
IYinaMzv1SexOjZq14OvWPgvz6WWjPanAckL//lNcLM+ejtN2KX5gJRtearEFZJsP+CmkfkjDtAP
o/05yv8BDT9BAapEZJtsINstAiiHBLxLaL9+e0XXnlwcu4X2LOFBZJIz+SjtrowLfmwDfyVmdXy/
OrXg4W2X2JsOaPke2vhMqOAvqvbfkk92hgSI2DHMYTsJTbtsW0dqzpgzzjbHBVT9To1VPvHhV83W
YtjSXUxeaGJMh0C6GXE/DDXYxpmZHUmkt/BLCZ4GMeImv5nl8G1vmgKj5WfjMo77kIYQv5W49R11
/e3usQrJ3kupD4D32NRID87gzrZXSUQhxkX1TDwCV3yW5g2FKsrkO8hTU4+39JB9fsvAnbDZdq8L
aTNJ0XUO5Li7tE/qyyuO6GK3ZIrCaR1nqQIHQ2ygIi2GWgyu0RsSSdQZ35SZZhOLukjYQ6T/8P88
nhz+KTx0QHXeKTvDLEWyOBBib6yhGVrmksbQiUadUtgPxchIPrAGi2N2F0tSAwWbwuqy1i3Dirz2
S8LZJ+gW+ZRsvyTbarHBewEbT6YbqVPAYuOkLYCCnh3JQYni7/TimowwsrM6R959LohfAy4wzU6R
GAiNetUaP2W5w/OjoIJzobRVV0KZa0zQxpIDBM1oJcgVHjqn3nsFQrFJGC0EEFCV7JBD3ukJiYpZ
x4vtJfhsASa79TGORSTArZMFV4nph8mYsvVOmFsXBx7eaJC3sSCaVLVZ32Qc647kfdE71SduiGPP
tkKBQE99v/ND4fxnOi272ejeiOMz+iDYTl0jn/rPFtCQuOA7AccRcNBE0decL5mwsuJSD4kdittc
YnmojLyCKGQhgLPJBJ2pLP29zRl6/YW11B3tlzt2m8PCFWZv2Ey51yxzjpwLhSm9WwsGf5FAdt3h
AnxTmmhngdj6oeUdUQ0kwj/ccTielsHcagSIcueGzk1/kkhx+sKZ5MWA50G4AWRv463pzduZsN7+
tqZHPL81dfipF2QFFC044afC+uGm/3a2XOGvPi2kMt2iAdiDZdGYyKPsHhErPxfleq5vZyiqeJb3
6vf+zj3Y9BWUuYLxZPYai7tQWBuYYVVs72DiUsXuIcG3dT6eu/HmNgmmjhnJaoKJFOr8zEQrKMMr
2qBwL7m4DdORE2Qk/hxkWIgeTrf+IEa3D+JNBy1aem3hlL4gLtqXWlalymziPTj1YDEwrgWpbkAx
9he27bJQ0/N1YKd2pERAnFrQUsioxcOVIub1AZ8NxeHRZ7kQf6hALcPI+M8yJjfjnwRXxTj+6sGb
cBW4zsinFrC0QINqHWp1AsaYQs3IIDhlXPmWupakTBLmcyIVsKlWhJ+HNl8iGjyGyNjJ06ytK325
ABW8hUgkuGc/sopHK5CxJy4ccdpKLfMPOHugJLvnbvr7mT8wqHysuAJ6PMbdSjgOQzv78ev3sRlw
NwAmlpnCfnD8/37Xbg6tnEbrEzokvgm32Oi1Nzq5f8AcNjwxYR0SBoHArCbjF5WYVHBLVXXJJF5E
zesGlJlXfexQyZLIVfqffGzGXUBWsNCoBlOVJ4hugpCnAVRUZNbD8OIBjtAkmpxn7q7dlSXNWXrb
QrahGbfZJUJId5PqOWtXYguPO3e4yV03OQolpuHO6T4Cb1WLLrmSzTXzp9DxL8RTWGyF+n/PYvmM
mnhy5/zMQhXxgXUIlKizhP2BWoP5HS1gzy6xWr/MR4DF6NPtz/d1I0S/B0ZOLsWROLsGq7TtrC9h
DweHtL4sC8RR4dFqrDzi+dGuioz5+bGJgXVDorFM6BIRZsVZoD3FcPZMkfmAY3IjPpnyNsDdGjFn
dOL0Cfc+RguUyHd1sKO/j/+xkfCQ/M2CYA+Al/iCFficAi7tFvvC7nWdQppK/Ik8wWm3rqjd79gX
BSqIoR3QWwP+1YCKzqZIBMJ1nvoNOfMuPAZSvux2E7ElK6Pvhp+4TFb0bkOkSVH8KY75/U08Uczv
iK5BOGz5sDYq/zsQnHAOcMr2q9v9r/obZlr+q21Yqd82tY/C8qUYdnpirIw/YxZ/FksaNc0ikLaj
rxAe+3urJ7qK273eRBoii0zHZ+Ym44qxBR9w1KlPawihkEr0LQDim9E1E4CH+57dtTSRrJZCJSZK
DApgERHhQMw0NTL5XijjXVWfBRBGqyLIq+PKbJszknOaMzISN3j6LMNk6jQ8hCafR5SWHjLQBE4n
M/FDSZTZmxfexvhFmPb+J2dEMdX+sRhCojjZTNS/m1/5PBPzQJgtE646CpyRNX/F0eMI/49Dm8XU
J9IFDD43AoFu8Umoq6G+W/beuQNhaHQt4Z/kgD/E0F1kKcymHLNxF70IgW3VT+UbxZpHuj5dLxcU
kzQILXel76r7ayZSjBVgJl5YxB7gI6GJG7e11s+tAZvaL6pQFvaP8T4cuGphe51lg2nRHSSR0IaQ
au56IWqlf0OhCEwncWTj+tTgVCUtRv2NQTh/3vLaFW43tf7AB+TT1UJ325C791alnQw8hb3XOlyU
zvNPU84IJ0vcHbd29zhyG/zEeAKUXi1pl0h/0PpP9MzMnAVXnXNuk9deDH+UZQKR3+CCkCSHUpHW
ld0Ju4+nApY2JQTgBeeif0onz6ISdTjMjAgSZj14OxLuCVyNIKCClM827DsqlFsfUOhQh3FtvhQ2
M8ERAkpRiytHYYcxrpRM/m5rnQxE7GA/Hf5nsJMIWEeloqWTJSZEj8APY5O3SyoWPO+ZtM3pDwg9
1AVAG5ah1/Vx43Cek+iR6YtShdN/HTLZxlBuoO3AU4qPRjI634XOlfEruK32bSOrte++YgtIXH0L
N5+4qY6Dh++8hhMxULS8MujbJSOcCmPr5TR7phzNbNnVHbHLpSvA+xXhBg2zue+3NtSWiYq28msR
xyDTVzNLGhY03+wJxLa0N1PqnlNdaIepA8bTlxxWh95VCGi8joy5z4r/HCg6S2sYYRLLKO27uvUw
vjSD6yd/eYLfPsfUFzlJo0WHqDdiXuF/0t2eu9AKm4Knj0jiTO/fJO25/4xv+9IpxCqdQxRrez0D
f4UXtgkF/zc0e1tjyqB+dPKQHZdjY1imaS/YSUriKH3mQRsDOhxnDbJTAmO8/P3gSU1XVNNj6nBh
ighZB+pSQ94WikTNPHiWEBo7m8LxWyJgZ0zQgXZr9QfjlBYiWdK7HLDSyJvUP9pujKnpQ2mB4fOH
HoZ3ofP1mcZrS5GzZ+daioqA8fWR1ym1eEHroQkcSY+0NzHlS0OfJgNkJGcm8gUKsleLv4lXzwIc
khq0h+qZXFDe4FEGOKrsox5FfLMFoE+Rtn5IRzWbGFwG0khlopm4mGsWgq2PgwfF0F55NHPdM6tr
T6G33LjCaETRSSPrZ++JsrAURKMdYCLYV1xbJpF6VzTuB2Jh2/SwJ5IRHp0tHGBd0o3yTjTmCdCP
+Bq0Woh9vqqO6+vi6r9RS+ysvo0prRq4THvOAegzbOlq+m2IDvCAHR2uynOFoASxvFRfjveZMbqn
c4sKgFdBiAgECV+Y6i5zN6+Yqe223vERMAu4K6AKdO9MH8nEUHQv1bhniyvexOTxaSbEMaR2devc
vH/G561gjSt/LLp7Zu/vxmEiM5JTw9K6HdV8FpzEHRj/zhqautkp+eoS3aTVNLca8fl2hFtp/oQ4
LfGcGekmszjHXViwiI7REFhGFr4NcLvt8ZW7Czxk4OnvO3huIHEClp+O9zmTWENesv0TnRCS9QJB
hdySLMUrLB1DnaP5yNWTWoPPFGYQFtcDvIHUYRicohyfaSXov4qLXuWsDXGYPOacYHwdp5hjAjUt
e8DRZSdu5KrGe4VamSKLf/1JYyA4OLLTvprP54RiGjA+/w8pnR5Kcib0FMuoKmsCS2IxsrZl2DWP
OGNa5mLdSGQ6kN7VnG1+e3nTB+fOgRusub3L0GfkCqdyWsXMJDDi5ulGFPJ2EKAKXXyt3QEp5J5+
fuKIdOeEiXzfPYekGPsapi5y8oebcPb3UGPwEZhQnuI9mgSXO4yewJrGCdEf/pkp4NTUjMU39Y6d
6JJ6FRcC/agLnu4Lp5utPppO+ilJvJCoTOdmPB1p18NCbkCETvyveCVx4T3BEx44YI4kOJP+H8GB
OSI7QgNXnIxTtKQkUYXP3BUSnstL36amJDTkHbCsUpLWfhETz8uGK0u2DtoEOAm9mjtunLD69dW9
VPBNoypnJO9gX0vOdIploAZ9M3Zp7bmoe0u86KE9CZ5WufGffeQzmK4F+NH/kmltNKmxWg90gvQ4
kGNLjCSaRFex3vhpO1wn3cs+DH5Dva3WTUw/1NtuFYcZOcNExTzvZ3D2Nr9U0q1w8LnMM57IUelT
RuZBziXCbj8t7zUfRI1zBP/b3IvAfhJlxmOWHEtRwzLOsRy+S87dBQ7VxK/8ZUBoaCKBcNNwd4Xd
ZMac4UddpbJrv00BqXHImhhJ+vLwQtSdW2Kdu+r7qnZKty9mE2XPZYNzMw8bG5+Z35xr1HaIfNgc
dBMgCLkRX0cC8PRnpbqRvaSYT7T0tbtN+YPZaM4nlgA4Nqbkupgskc7hg8TNTVESMG/GQU8fV3kN
KTQ7QmV+crfeBXpic26mU3v7LXsCGyuoV4sVSwaZn9/AVMnfmTEILpJfiKbjZH0jD0Z089KcKQKi
fYMz/qNDHGVo/RsJuA9v9T+1DwFQTNnWD1hNxCBgEIJ580GPzim1Uc9FORa6juNQ44aXe7PC2KzJ
W0yQpbAqjUj/v+HzTCW7kbYYBUSV6FG8a9/IAOBFvbDBNDkKxqSI+MzW7VdM0RBhprfXP6szRzi7
TYxKYpuJCLsyG62EF5xI/UC3BwcR6OLzWqQdHMfyUMoCDuL9bQSS0amZue5CbOSO9yz/GCyNCH5/
OnC1uar/RrwXwjGby9LmYOxbl5oGN/Ob/wcamEZ46lORaQaGt+uzx7JW8rYcfDIEL/OF3qJqfjA9
yZNdIaggGJIUu8tFQ3Pe+SdQti7JBFpDOm+IA2K6iIFcX3hwB29wnQaMN3BAMOANPs/OiFt9sSdR
/rulRCv3IfQXLdBesjcVBiMO0ZC555HJfRYPLY7gGvq2AKra8yqstw9TYfDmACbQJt5xcc0/QAeI
9iUdLf0imlbMjDf9OWsqa2BOvwIEAdXQwvaumWYx3LKSWK/Gtlt3bQPIemtq43/BYgiGsjhssR3f
ANhSSsc+8UCfnoUlOPEalHMCNtAUBdvDfPQhl71tTsEYFU7VtvjaMvG2N4F8s88xyw05eMzHbflC
m9rVf/ywfJ19XwFTebLTxSlKbAmq8s4uYbHEo8uh2suICOTmhpbTVZ9vAzGrMoWry/dAvcO3r4im
PiVuzMYWWHybxnZCadKIlPwEMXMFK1zSy7mqBMsMOExLwim81CL1vtMjXVj5LqBazo1bKjkj9BUf
GZTyulUW6H2WCBq4eQcf3JdgO+0cp3+dBe4nCyq7vQk3oylryUgLTVZnB4fQlLlmJFuDmdyFYRZk
0jzC5Xjv29RQYzN/Ob43K6c04oyU4EFxq927bBWl7UWO3LoT1CxxeUCvGKpHZRw8qRRxffFoWc8N
ZA244Y1b+KxYD5XhiIKgcdNrNEs1h+MbXR7pb3MI8LdcxXgiHUCpA19ZGjoS1w4Luyu5xJqs5l7a
EtJ5xQ0cw4njb1nfkxKv3sKsHa0yqO2ZiSnSbN6jgkWpnFr1NIuOyXLa3QBgyd0C6T1wGhYlFfHQ
pXXyls60DP8xEoDzWHGyCBArrn3kuu+zB/SbBVvSR3dHWNQM6pkZatKn7MZfY6Re8G4t1HOJ87kZ
otP32HcQNIU03w7n4z7O+rCTRda+oku85a+mHY2O//eSKz4Mt/hvACPMVWjTK5BZagKK7aPs6vdf
HWdPcz/ltt/HFE8Y+VeNSauQ7RiHimMAXjFGm9RsW2V/dHLokH9F+f5iOnjpDzwNoNsVbGDeS7sQ
pjQovimrGtlclwso2psBRWv5bsuKEG3wU3/3EFEaeHcnZHqyGst04pzNkbGT9m5bHyLAOdL9yjuC
zs9xIhaon9U4VkE08NWbpMbA4wpeyd6cQt7Slm/xJetJ66K1hdormXD/Htz02CXxc5FRkrB0HC5O
yimi3J7GPv6rw4Lwkhxo/ZgS1T1lhEwIi52XxFe3CjEtTZuJij6Ylkz2PusHjh8Axz5rWHkTcp/V
EQYY4L4IbBGKqlxf7+Gf68djHjBBjczoO8mh3K1l5GqgH/+y1R4L+0s2D1EB9nruMc1IgntBCzjB
yVnG6kTJ8f+7Mh4eRntGdY1a27ttX/tAArztQq7h5c1hM3KqZc2xE6J51WKGDZDetFfIf1pdstSd
zo/X3MU8ZNdpYf+YOQ62F7lkg/fd0ifNyZyjl8CT1hlLXpBObxWa3KbntNqxxP6cWYcigRiqnxy+
GMF4iUZxbTGbze4ZzJobxPcHFrvDyrrlfIsuV7SKrDRvbpQgChJDp+g0i/Bcolx3cvuTh7H2Q9Yn
C4pL14aG0cm6HIcwQ2oIVdum4poubPW0uIUVUpXQBwipD4q5P5MOCE6wi5WGniprVPcY/2F7IzEI
yR7FGEdtdcFkS58VpjkDsQPO3MbWVWHcHOwgjgin0k4JTGBKyX5IWo1sHj17eizbk42zZ/vEJLpj
IR/oWyg5pAJDvHx6pgXKRgry+Ejs4Jtzq67hAsQ/ldpbblGQPQQTk1ww+eyHSMSoK5g0AouwUC6l
L4+MWMRfxlVSE0LNuoKrJYGjVOPwM45efUeMIIdNAWMR0b+IbtrmCam164kZIvRQLRGAgL/+NDXR
fA6LGN4bdNoaqJ1Ud1HXLX9wr2MIsT5sS3bNk7NuWaXey+wt3dsrP8UEnuhgppjFHmel/DoE3mgy
usc+Ud1Wa5rFcRHEqfbk23Df5vV6E2qoP3y+GqTzAsdib1OZyuHWCLOY6GGaAkdLaP1d5EDn0dY+
fEhxEnabl2YrnrfI/YeRvlRSh738CrLbgVaZzOT0ptAQ9G+JLcG4v5cVOBBbddB9OeDiK+JN18FI
KRBMnvvLRDSORmdjHN8XFG4Hug29dDV7Y9ke8tbv9efUaXBr92EEWVYuBxXEiIaCqfSHni2TAYe+
pl4JxDg6YxOI7j8NokV9gPI09tAS8I8h/LOIqXkpO71kLBaMiob5f8U8qq3UgnwkVPR7ldNQQSJp
qMuQu6r4MPR8LpU3fzCTvRJoEOFAh8JhTHc073anK1m9SgZgcAk2OHUXXtoQfJ5ptpmDE3pw9tiq
133KFO9pAiZvYmFKaMbulAdziMXo+BhTOIpcg5OkENiq3etbzs7XQcpulcDhoq81YomGw+XqJEJA
3q2/Jc2JlzIiBLeu/4w0Z676m2aw0F6/TPCOCPIzrURAx6mGmnWANynBQVw8rkr3RxjnAYuZ+3qd
YbTGKp1EBI7t+z2ZLf4z+qg5LVL1x+74lcs86OiwFj0DQFEhfd3INRbhNZQtlEZpApg70Ivc7HnR
AWAn2zBhP9MfnivgI3qHWGXiOZBM2fWPraFIY+OHy/A9+qaoFpH5qYTe8xKOQdQl37jCHNjJNWk1
jbPgySN77KPXBiZ2Ip6zQTIb/mNv4V0Kw2kTHfB3hMZU8junrgFXuCHO5H3WozTc3/jeOYWdzEKR
PxXJcAULYTPY6eEO6xNqsY9XKCI0hMGoJmp+hDq+7bxeJDjh13I1XEcsFiqIQLZuk2y06qjeYa07
nyApVw7HOdUhjXEOJ25juIZvzybWLDZ8aBbbHEKTt1XrYA3HdNykQr/MP7Nap/WARsdlNOas3vkt
VLIedjlCsmcdHRtoKOO4qqyBuO2MqLtJv/kVHBXB1nbYkLUccTG6+vTe5qW/UBCSateOn3om20V8
sH3Om+CDu9v4xftPhVeshKaPYFrUgDGVQwAPOgGWlbDoCVho1IWZDWcbV5Tj4HDX9297sU0zW/8V
QIGahJgYwWYQcx5vMBI0oUWt2+rrdBWB7gRHLFiCuSO6vAlh7Y3+7y8KAgS/9FJJbtKzhtdvoecb
c8aWVZmDM35ChWogK2mfeTab/XbSPJatzgSbZEHdVxgmUOi8ShHjYnAakLvaVKiEcf/ULPGVtQh2
SdGs317CKSDG4+fRmnJpzjAFobWUddWIdgc9tDhRLFEyyRPKHPeEQvw/dguvmNsgvDDbfZCdfcvf
qX9KjyY0Cj9iHCeIDpMvsGjiLv2Wo+d50LwoNOWZtfCw1pWj5Qu8L9dU89t7Gi99Dnwxv1WL/QYt
BH0pnNOmZHScOuQTzZbJEGjwVnko7tMwQ40L2vqYyiEP2e2sCP3akCcHzMuigrwaQvicithjqc9o
1iH/FPvVjezHHWO7+nQj5YNII9WH5+kiXC06YoQMtdYGuTHI8f4n9DFKADInLHZv3fvRcHrlHRhv
tYP35D3Gg1a4S4mPsCx6NexeNITPiKKMEl2hq4/IcaOImJUbY8ymAOLhut0cz7wLEebdLn390Bbc
vgl4bwSgBLQsshGhy0UkbA13B9v8PGRZIYmVVMBoFT8ZgpIXPNBu7pLhsKu4Z5QCDgH30rWR+jri
bT/N8VCUp2de70iPmdujt8bohGzt0hgRsoQJf7Fc2hqdidqsjeUMuNYKJQmRX0e0YRxa6lyF2RrF
bsU8eXrwx1CUvtY7CSKgPe2YAE60zoq9Vp96V8MowU6rRueCLd83x4KVsulHZqcnFR7Qj2Eqfvod
ttCNbAu8NNg+nrxNdgv1pbmqv3xqc5Tn6XWD2Yg8GKx53bdySAjjhT5hLVAiFGv7UwYZzo2tOkvH
YRZs7ekVRvOwKN3vkMlNfCgVkAeD/P7Fa5zBbeWzTvWQGkEFFyw/yRGAHOfSwHjiMLT8bjFb9AUP
+mNuoNS5VEBjACISQ5czgJniFhj4cYVZpjsXCtGzWTn4F11Cw53deZPTxnlcVBIceaWHKW72gajQ
cKgGFBzDkSIBmYN8pcxM4691e3zgqPrvp9eZhdMcGp8vRgOTCHoSYPA0Bk+IvazsUcFNOABeKm7E
T+ceK9lvZTfBIEZaxuxMljDL7H3Ip4YzPOJlD5QJhiPT/AGpA9J3rJRLuwGVNrOk7DuSpernptsA
pmVsfJKRXDf23D/nVtmF9cSO9hkKsdTxl5LiI6ALmV8WZ7Gif2gRh05nAnEfCmzAqDZd/+RQ8AOn
X1h5zxnYuGCIB86tCL7JctysCKd1b/Md65DxFSGPvUcEsyeaPKd7S364GVZ8kQwRzX5j9zZKPHam
F/8hdsAnQGkcgXnz3cUXqPLLu7jSUbUES60kNUNP11pZibkOr2zRvVyYspkCjyHsv5EY3fi5XM3+
lgwsvMRsw37b+Kq0tTv+S2WQDgSWus1cfzrri3qKJK6YOkpS+sHXSsM8sLj1+sd0LXYxrOV4gVxb
1rXUhVf+4jyXrxBIThq34bIbtUsQ2uKV40BSPahgHDtffsXVbzNgKeIZQ0xP7kSAAtbDl5toThXB
Sf3CgEK410uef0Q82tP4pzxafYu/oBLblaYuLJdUYp9xNkj9mv53OSZwT4gThJ2KBt5YEy+wGy2l
Dy1CEpRdKgEf7vwlHS82mG2xG7FSminFMv8JMVkOIOdjCd0+obR1P4gUN48IVqC1/yapSQZJ5GZA
MJBKVLV9wg/oIGAyHLwuqiG68s+Edg/vBvaTCBYO+nDzwu+aH2dHF0LbazafSFy+ZJNVkpGfwYkO
DHhAaF7xvVmm+2Uh5qvVkG3BQAk/tcqcHvg+kUlrK0EpwmYHKbOpGRhglf06nHWalnm2kJEuMR0H
Zx1Gt60ur/f5bFjBTrvD8n9d02KczfY0u1vmlWQKfNaXkJ3QPZfew87ecfbyT7yiQy5UxPcsPpmK
BAOMdXkC02cOr4dH8+vUGLo6DwZfp1LwVUellPZI2mYp1HBuz1DSIQ3LLFrV1J+iJtufRJsNO7zl
u3fFexnEyyIxXPfvRBtmYlT2uOFj9FfCRO2NwGvpMsugnpKfn6ASjouu/L728OdZF4WYK1CpPfE+
bORNcw2QUnnDlK8QthR5n/Cue00jlmi1a+AG5E5LUXm5XoZh44fXskPsLLbOIvY4/Sd6mjF0YSC2
4/In01vVx1SW4tslVVNlll5uMpcCUhwTblcWMFQAkDOxXGL9CX8H+8oG+t38ZO+UxonaUXmoiJAm
q8S3WrJdRUuHUwccig7OQ5xlMlAHoCFGcmaVa9DsZGAFk9XJvi9nUVFoqKcBxrJpybUN7nt58OOJ
vKz4Kmr/67BtbqMQyHQiqiVfftyv2JhqAJqBF9/rGsm6IA1GFGexnj7JRd/X4QQQRvpQU4nSdjcg
j7/Q/PeAF+jx8/ZscDbPx6/0yp9BK57jdQpsrRpGx90YCWPuA2BTl9QkbCTDnMIKCvKbjlKjBiry
mX04oE+i56nZ/zLgPnTk+DM70UqH7dddEAUYaCmwIyoYDzzNupQAlSmQgDsG0zFyLgipWwdiL99E
Jkqa3YKaOZ5zHtj2UfZCSOHiwRzZzP0DbU51vu/Mfn8LKwCf2zg2MreSxQ4JsHbovX7QWOBR9ML1
5BxnO/gFATZI8zKIm2bF0VN+2AjILMLK5wL+zIHO4D/+3HCGl7ptsl+Tt5E1vbeE9XM9qBxxrSx6
UYvgadEc7kWuapiQ/SYfuo7S8nAOjwskvVgLavGsOGmwa5OwDkoAl/LttqZqoYFpLkqXs/26+w1k
JsxHf0SsipaDqQBtffOZ3nFyvJhcYZTR3jBQuRL2+/o+Jjy1J8QQBrTPWNhvsk8NKBC4lZx1+pjP
/z76uWqjYOgSTpDAYyFDwZt9OCzovKALiRSWYr2rIQ9TzZnHBf7/VxfN6XPO4I270Hvf5CG1WDKu
hs/JQQhxWKuvXcsgziEts10UeDiDBkEo2JbPXPloGp2RgeWK5q6XixmHG8iH+EDHSo4lia7XmRlT
72N+V3vbr2VyJRsIjnA2558DnLj97mb31la6nshhosj+Ib51WgaGvGgLsDj4FJLOJpAp2iZ8w/gf
bSnVbi8HygoJ+O+5A5DzOomYUnG43qRKQyz++WNU5Inqs3qp1pjpFX5KuyNUf6/bHev/yPG1OK5x
anuCXjnpcuUXuMT/AaFp10UvcK8eExWSxeWV/CNlZ9Imy2DRcqDBxj8XiuuJBwW8ZkWg0BTIfIH+
bG0nu+klsbN2EKpkNdXQ5FeRZKf3+0ldowRoOIAQvJ0DkPs859H+yYeeNWl18mghGKq2S8eixfEZ
FTHAXnDVfFr1X7rr2RLsp+TQ/5dudjhxrxikmVuyLstK6GVBEtjCvSThwpNMewFmw6VGw1hu69Jy
eqg6SFIn0sJcioYMgpgOP8PlJT6RYx7Mvw06un3pYM6jIEFTH4aUB7obtvNdJkjc6A37Qbi5W0SO
tPgtrh56/Y/8/fK5KH6UnC5MWuwaQh91C6wAQgELT2nO8/moBWUhtSWId/nOylRMGJPnZuTjCEoi
wYBmSby68+x2ZpY8WbFKGbjC0gG0OP34pXv86x1x0YxWxhSnvzGs9qA3yo32gvYCykyMwV8AqiW6
0Dipc7Xslccs9vq7yEic4OD+AGlMgQbW3W+QQ6PnNZcmM9eYstZdl4rlh7QObebyjYYVRsjOStLd
BqeexMjd27liJ9K2FLK84eLAYLCfQ7s+epKgdvx5dLTDZyYFsXgfaRE96heaPzRcurQOTcRVe00b
O9Ko2Gb69+lyuRP/aUcV5g4cH6rUhYdNcnrQMYx4FIBXkjpP8VgrG4G0ncofmjfsuMVn1OLfZKHa
RVJUCyFNim7Zxijv0ccGSGZT48ruq8Ft/IDdfnU2yBpH9YqOyoKv2jfRoUO1NPiabizo5b5MMyPh
j7rDQ/0zEGrmy7inxg3sapWgT8AE8JkBrVdAXbRY46/8P2rwax8m6dYHs9vheeOBq7Wi/ne2vbMG
CqCwNP7vAgoe51xYycw0ouQRRM4+Bg4SYXOW5oKpHpYgGNGIUjAJnTrBUFJfS7QobK2/n/OKsxwn
BVJ+dWfAKM0lW/SofIMY7CAE1jGsppe1XHWFxU4dClD6VW5JB38YR+kmzn1G6HBieKxleit5w5So
3EH37V3KCyuWjNyXHSrfUqFzy3o5IdRJg55tR3GQfK3AlvuOSuDnzTL0RXavmaqhZrRqAniJg866
hS84h0sbJ2OpORcXv3hTM8Oa3FvkRihRmk4OOOaLmjNw5AFJ82Kw3aWwGBP/XBTFhkLo++aI6rpO
WPykkqCE1bjewPsQL7rYSJIRnqk4nckt4Ed0yeOBp+S1caJlNMew/E6eVucvylFFA0sKy2G6APwX
rVGOV7HUHjblPYcRUbvhIgZ3SorVLTzIby+qNypSUILOxzdjiKm0iH4OkZ873C/tnntstRx9VzRE
cZ6bRYT2h4D/R3YjaMF2upNDRGpP4yM3cqW4tFQ3q8fkkYY05Nv3h7PKBvp9p+mMvKU/SJEqjpmc
NdELEX8qeRqLBXEj7+gHChqzHC6Jy/rRtGQTmoe4Efw6QJ+icMFbPLgb/ds8M43DQzavTpQYSysa
L/oHsThP8kvgXXcUlp5sSnvSzyjlUIs9yQUceJXDd6kktw3CqEixinadsmTUf9RrePMRIXlZf6uP
8+zClL7fNour566Msyta4V6sa33HjZxLjhuHR/y+5CcLdJSkjYwm4SVLisieAJkgbP5ugKXzQMJy
p+oBmnVVddR1mtrfjisgTguC8Yw/iY8kXJtjRJa8zrhWDJQtTfSlDk3Mbafa3JrvJMwHGMHFbtZ/
Ddf2sN8lN5nRvUTtIOx3HvwtyzuLeoM4hCkaonmnXkzzNiwg+/SaeFpRcFY22eV1hOm40XqnTl6v
Ch+peCOQPeGW+gPv9MHcGWOfhRzjkvqypQCS7tjROIX9O4smG0Tb8OgMLBFtRjzkYPj7mD0mHURq
Elj8Hx7kopMXb+g/nR+uBE1icmQgfvMKnY0a5cFb/OXrm09lO1jD/BSJBWGGaqpeRAFos3EWsYUD
AyshKKaSv3vkv9ZlqkM7ylAfmZe9c0k1JqnMr/1uYa1cptPrKzF+Z2SNx45HlFi/5itw3FDkZTQ4
9F7d9gicOFv4sk91GtY4u87ji1fPz4CyiHLF6ygJRWLNhb9Ooh0PHABVE1DVGyDuFCTB5ibTSP6Z
lpijMtXogvtHkefCP275AvXsrhQbtSnUUmfXoUP+NEIgz8cwloHAj4Rjx8dTHquG0WQSpDrmcrI3
bAfXMW/+B930KhTyD55L+86EhbUYbqokI8EfbQZ8mJ7a/H4QFWBhunW5SupxYf2uRxRNycwf5Rv6
nN5gmxEYh8ZJkXYXBF+VccTFnRMpz5Fg34Mhlv2pnFt4DX+/Scy0PPVE2gTFjMgyefHJC3m8XZKW
pU7NvfoNwavXsaR/RtLJsfsSTX6qhE2Yv+u3VxE/vRN2FYCNOoNUl1EErkwjmQrtk9lrEStsO0Tt
HfNh/uSzFRBSI8n5PXL8sGGH6Na2xHbrjpmsy/Aai9bw3/cX4v5Qldj8jIm3SX3R3tqXaFHa2JIt
4rmbmoDbKkZ3ln6jDIb1FjFvMk4Xk1wHQRlc5r/LQD6VxsI1FNbo5e8dwUK7CyHFYRatEvP1Ae7q
KGavgXvYCwD5T2zP2ACS7trcXadmSuuY1UFalKOUOJbHr3UodZAIPP8YhlrGcX2C7qvy7t+z8BRa
qNjbwaNENOpusc0j5Wa5Rs/jDzxb+VjSN/M/B8BegX8yS5ZN8+H8gd4V1VVCg7h1P98ab+Hs3RE+
1tcDrapGzQk2ps2ULFLDnjlCJ0vBk3CslylTN7FICUHRdSydzYoL9eacMyTKNz/ruW2SISHLPp21
j3kfJUuimrmW2dgFysd+JZfdE5BCKGDGtBEgr3Pp/mLVC2y1UsAs003FqHjhw56XkHY7jaIVLrSC
S6NL6ms0enbm59+PvZVo8STUzoLpUiLIj4nB9jn1l7gyqf6Edl4C/BxIVJfrdxiyHz+NYT05GdF7
t0pR0Tc2NzL0cJ+ZpMXR6SwJBiNFPAEzDa4CEcnnY8oaZ42WF4MI2hcg0k5pqwzgdtbILETNJHNH
7XMmeZBIINATYzQbmQRZvr9A9A1AvvVKD+S3/yCqryMzQ9opno28kmHUFMouzFy7xxe2u7ztK3yl
9o8QbofkZAbxI6Ez4QPYp7YQyqYVDF/4tWe9l1MMfZsG2wdVadSVURDn2RLmtEAA9H4b+PshWam3
p0fCfJwOGwSajlds3i09KWpa9MuuH4UMVkhd00L05lZNYQIGbrDcPjkR7pNt8a3ElFWwlQQwDr3x
7BS6ezRQa0Gl5rD33D79aOK7owGj0XxWQYzB2k+6W8cMiFR1Ls8ZKXV1hKbsa0dPGayTNXeqA2Rt
jIXq3tmylVP1+W0BWDOKn6WDa4283wNV2nkW0uFKbN8Xp9BtVWRC044q5z4/QcV95xgGCp0Zht1X
59kzZXqbLSFZg9y4aBjD4+hnMjryrnC4WY/vXm3FvYmmUFSDZUrQsgZaoZufyD3WXgmAGArBn4Gc
KvXzSBQ2qj8VM/q1lu+YPoTR3xHr6qYPbxV7DRNgUS5e8pPDbOEAXXX9zSMfJImcDiabWg4VT5HO
UP2JyEoEfkeXdKET+Wm1Oi9AjLgAHuv4EcAimSqTfq0NVOAveAnYcyJEqb2WUJeUCLf9rvjy8tAw
9FxVYZM+uVt4WG/Q9iBvFhUr4Nw8xtC8hpuV4RfaaxXur24m609EALp/AAn7K+pOFiqDy71k+i3X
/vr9ILw/2vsc5Cn2+e+g5Wq2G3r5F1MCZ4gcth02SgOcucGYT2HBlFEXnE5tYGePqzwxnDyH7Nd3
WhBYkD0ej+kue8OO3335mDq0/W9Xpk5Mvja7Kw8Etn8kdm0ComQz1CG15/G3gN0pTKtJPZSbkBAU
HaHmNFnUg99Dgwnv9bMIIcQpyUxuCmZHmglvOmP8QCeEd5+xhcJj04LZFdsoNhLCoYUPrw14cNu6
vFBQFaZ0q5NCmIoKrbQxH9aNl5k3FGjT3UGniHGWTm2F+CE40hQk3k9NCyANK4YQv1DAeHYmFSeL
pzOLkYAlBprDdo4RzmeSFzbbQfrLiiO0HSFpxwp82LIAPr3970qr9teJiIsT1pKspI79DRj/oIHJ
oTlFQ56tTCipeMFW5XeprXdV6xouyzBYCc5agyc7YRuczD5wSx0wLkH0Dy/RdWH74tFlIbQmwwdI
BKw/v9+Z+GBmeOWCYIm6pPRHXyTaMPrF6Hrq8C6pa+1/w9hsbRSbY20impcYZ8BChuqKpe6M91vo
enDPpKBdOccRmEsu9DMhIbVVzp3nYFYHof3z9m+bX3JcsdL1H1wPHTBlBNHPoXrJTSm6J6N73gsC
w4J+fqejd7OwtwgalayKhWEI7YClT0Wko5ni0DIloFQnowgAfi++x9TC2KbbMj7esvI1kUkUQcQ5
SJhNqGZJON8BTcnQVk5Sv8FFbZrYrCjRXBfSXG3WxXCLT2d1Z1dr0gFzBMN1VeK4BNd9Ur8bZEoZ
ZiL0B/QhmLaLt1pxg/PqEXv/Ztl8VI5M2vOvKVAIearWcumn2wQ+kcqo+4IDy1rY41YaVrS9FABA
Pi1pieYoC1f4Z9BrCa89IuHkpu/9QbcxLn3iN6lwnOwZNHUIPTXZzDA2gXefbPIFI+baHARqbtdp
b2/gcAYc5m8ihLptgU1ciE1MZeqmWDTFn3iXVV8mlJLha7bD8NyYsKPdtriSZXiwKJwUr1dfPg08
/JCQ7yIrwTSqdSPT7x4Ex6UraDlthF3edrmzy3nt12GUOQ5PrhCBqbGzTxKVpeHF+Gty3kSjuF5g
4MIJVWmd1NP08yr2KU/rfAK9q9G/YccvB2o9i1dvAxp3iU+3/+0WN5VyCzo2TCGVyCBmE/WaQav1
zTXX9I6ax/ASbltggYqdk00FeZlQXzLDHMHL8avzc2iK/933fiHNIfEfxOotpAG83kI1eD70BNKr
kCUsgYv3li8n4oLz+P9+uIM2O6zvbJ7bAwlbGcVWeHCyJSqd0MvHH67JEjfRYBtg5ZdiG0IwyCSb
Vivyj4k0VyZWOSPW2i5o1o9oB2mthonQddzIpN97bOMuaL/ppJeftJStKnfc+x2/rfhoqb5JOQKI
7K5MtP+MjujtXj6dffrN7A6d/udtw5WK4qQwbBPjFFxUh4U+I0ZU1Fmsz+cnF/2Yq7lfmhrPRUot
u8x/7PFhiqlSJY4TXzjIYLBuD5w+Bq1eEZfihNN9RcSLtgzymS8MwsHwZ655/I2WmBo8d42rqTho
WbrP3GIhWYN9DLmB1SslHjGs6V687eEUAmpQ2aXqnpBgOJu5xHGalPzEIze5JtjxQlO9+cbOX/wZ
KEw5zgEXzb7CdTdt1smy8BNTEGhRD4Hs3lUogu6ma10dTYu+oz3YlPDZbx+c/dd2r+A+kIqdwt9J
hZekL/BjobpdDdM++Dz7lj1jqDZFui/O8iCcrAAb4LvEZMUmYGvf0nmDnbDuouWij/YeINJmtNhl
KJ3vUR8DSNceGuzL7tiy1I3Q8w1jqSPFTWcAPKOz25YpbpsTGgNI0tr5kRkH9n0evzu5J72Rfe92
D4tfHwse1+WTyRc33xweGVTpISwk5tX5vUn7Lb/MmcNcF7yYwvqMhLuitCd5tuY6kotHog4O4TMo
nzirbGmfUDxn95xvz0qVs4sGE/JQ5DkC5SSlpHw0OYhL3HYj1RyEwTl3Miy9LDsVi+9RhnCmG0ct
nJzfHD+nYPtHo/R9k2Oas9MxEKDJ941EldmxAyDjkCwnIBasSQTYeAGqEE1BKR9GGNueEfbdpKF2
sBeBp78t4r6ToLf+sOOOF2SFTmCNqndqHZ7c7v20Q1E2gySk0XuF7egiXDVmJhqDcMHUnsGrHR/f
YPoDvhiyJh95fnZpxoI2bbwBrlU5B7JBqhRuMqQ5dX+sv5ca0aRfknbcrwB7v4aKPhqBX3x6zDs8
QmXowGx6V0bKpRg6k3jz3pSAH71DPalIYOz5zgQFB62f0L0SD4IEZf8kpy82TEwY4l+GR1cPl5Om
Wyx6EUyjNpU3jGfJflHm7OETgZIbpe5PZD01IOM6LqUvJHyzu0oIZvBvzG9+aqGYOqztQAQRDM8X
bd3xSqGYWhxBfv2KjIWZ/BF+qhOvrpmSP6xORGZaE0FLcwBeedPLqsvV0g/5AxvwQwx2le9bmWke
ggvwo3BW0BlsZc/BDiBMCsm4IcGtHdqnT+v+vv1Oji79eHW2A/XPJJnQV6sZzZN/MXhyHAAS8WX4
NTTKgLEM8yX36oei6K7IP3dU4qkvdggq7E2x0u9HkNoRQwqbQjlIlCqpeBSiov9doejBcjiIELia
XjOiUAOMHLIbEbONSdkjXZcZhqFtnTcWkMur311L8G3kilWnejIAhdM4Akm/VMEtm0qAwpUkhCfI
aHuK26hODJDeXexZddIUJhcA0FBizmJj/VYv/jLRb7o1pLCb+SL3xqrwXEf4VKMSDKeBaAlB8jVT
qGndR/uMNbDFzzJGFLo2dbd3FCTxObvSpUGrHkpv7PNr6M1UZwLWQGv4WYws5HjYVTzoeCNSm1dk
wPz95e69RKdmlM46HkR9CQJd2UydxWS2XdzdKxCwmXsxXlx4ZS1gLWa7MRPG/TCy0+xI9sOwWQ4h
wGqJK89lLbwygg88bW598pESlrLFfDbKg8f1vJyekRXr+cPsiEojaterc/8OtOGdX8X+riM3hsKE
9ooRoD8XCsOz1Vg1xhudNTtlKvhm+5KBe6Q1wxyxK+WH0v3CQxa7tmRhpywhQcx5Vdt49sb478VE
pTRnL6orK2E9CCph7ElB+BxkaDr487+hzKFZAB2XO711+ywCsloA1pQ42gpdlJI4aMHxTKjXOBtT
5hdTjS4TnQxcAWeSNmAjs75rdoX6Y4R0Tpu/91mc6pNtIWQfXSiaz+YM8DqSpileIULJnAGFHKsG
ongi2SxZs66+eP9UqavHqm16/SlHinxT/oezhOjdZX4eGYSmGYkz2yWHTOR9Lfw2+48D2IbK0k7l
fgdSXM6RQYHdxJeyEedSFZXgHB8giU0a9JxO1iiiuslqGe+kdqVPx5s+ja+JNjiF3PBJMKuvVerq
fMut8fG7PNe+T0gRJwJeosiCfat+5Wdt6OPagvI9vbz+cwpqUEX4Oc9cGkHmrdTr8JBiNs4JUpph
4W69qm/2QYaXyY9/8DYK8G6C/behl1Be4t9PtWToDs7bM6yPt/05u9dFlkftbC19haZ3cUgcinnP
Ul4sDr3UaLAfZ+ULN6L3hgiafMCw1+yGEaoZ7geN+x0EMdA5JEjx4ukdIlM2I0nJDVG9JyowK0zA
nFJx8lglqpRyw+h+gmc3rdadXcSi3g44YByqV5ze0f1L3rFrER2Jj7/vgLXn1AlCrIYXhjj87ctS
WIEWgh9W2KuHjSr+1Uj6F8su/bBVj0VKqyNOVxtsa3ePCqxad7i7XR/iqM7i1c/EiYXrn0Lv3MFU
QfLKrRNZVw0q5FTLvUZ60Fl+CkYBFtkK3UF9lXS19oeGpZz1kYymxMy/LQoQISzE+zSmD/yxWOUE
+N/9pcEqFZF4gtMp6HC+FSlbMw67zXjVzBWXZC2KqffTs8yMUQUa6eIFD2RzYCYSDwVE9acSM0CX
7djK4IUYHCuytNFidoo7ubGE2oDpSQOrcDiIzH85UzxM7mj5zn3ZNwJyvBUTw6ZczwR9BRDOyPnn
AMlreW2+xZCJroOuPImANPLSiabaAXeuagR/44KabXEMUjgWkvplGBTGOQ3ZOqFKMkEDOAErRDk4
RQ+uf9fQJP0zTN+iIPwYSHyQqyO0ddDEOjFEFDVP8bkXkBqJjiuke3WjTyL7+ur2ew1ui9Lta9Jn
+z4lwZjLT1+4ufbT/T0HYba6NHJcz+o8RDhW4L0+ogxQxL4oaUkuMumF15Vr4MsZg2DtCyvQlO9C
HiHKs/hCd9q4CnsrPR/AACTkj6z0HXbsBcM+/XEtMKgUyeD1Efn0nwdlOrjK1BPd+PwCi5Fqr8TP
b2hi3riIqmQWAb4vKny/nKqWWyeImYAzIHMZJI/MN9TBJ6RZCIpay4nUVUrrAvihaniPsYJH9SOu
sUTD1TMDrOPukjJLh9ttUY/+sYjcy2pEgheKgBHVQix5CQ3qQxSejNnkzKiTCDUrhoB8InaANiTi
+sekjgOX8gumTBg7wnGcDN5fKrYsSCi21muaj4NDJ0FVT1G8IIHHJ4ABaJAfoJnUhj0AEOgvYPGP
4v9DgS3AzlKRuL5hMgVYDLztfr1vxirOSJ5OkM1/ctcC46DiJkG0ubBVZF2i/vtWA2JhEuV8Xx5Z
yc8sg43bJdDWf/jCM0kGcTZK+RCDh6Js2tC88KnWtHVXWfNJfVovbpxOpRi554BhVi1LcUod3HNH
Pwp672C9k4KAzreAeKk/zltHF6ASuyJN1UfSWJD82UyddmV480dsDIfYNQ012+XMi3Q6jEzA56Kb
T60VPtZ3wPJ9HBAZnHqa4oxPUe7DvnLtSTZiqbL3Jf8aZzFnOncJ/AweSRbd19mvnHDBkAdyrzjW
1X3E8v4BtIV6jw1cgVlCJXvUaq9edVMEhp8DgA+zOFgjMPsTjmhUcz35a0sNeMLU9aRzuRMToJX5
capsH0CtYLzi/WALwjaYmb+ng9YBjQGPAIkef29pIly/xZiM9R8M5ovbuNQ0HpvDh9V5ZNVkKC4Y
ZuOIajJt9V15X8s/553DU9zCjH18w8gyEX0mKTU/yqZSO2TwJ3q7/z6uK2Op3YVL7cde7PSg0+Am
hf//5OAj6IpbIqcitoUFdjE4BIwzWTVJUYzkNBQY7sJA7nb22Fo+34lpVhhIte2+k3jRAMh1lQwy
5z34LwJCzuHmamYgfVG6HhkP2zavOYF6AssB6OGKyualgwkm6+7YpLm10g2njV0MLGj2PlQNhwAK
o8k1JAuXwshZ/oBN9cBd6bhiKmGUQuoEkIbQv11lUEV9HBF3i+129brWJAJTyulJvKv+UUJKz1e8
Ko5jzuy9FkmI2knIeGQg++lamYSbZh2zHKKzK/EX5ixfEmWyV7kjRmyFgH9QlN69VbhLvEox2Kbx
H7iS0M7gSsf7sAfmGSORyHYUAuiO8vNeWUi5l9M0RU+CFoN2VDWMXcydheuWouvl/Sgs4E4x60Xd
LRVXZR80qtGYxQVgVzdwmEIzu07fzv7aPIWzLXBrQ9IZiq6/Vb2ANCWoyFvr+4EDU2B9I8iW/QP5
+oUMM0fl7YBU/xw5arW9kTFEcEvzXgIt+AUq0BJKBe7wEiB7pHHFR3SrnVcCr0n67AagBQtIjDfO
yp/tg7vro8hgwJh5FhXUb5TNwrqYEzscMxPer915a2/I7sgya3L+SXmAe5Sk81hf+lMWVHKKCnvD
mvOMssE0YHnqhpiE40EuhlOqhgkvK20clPZTZfkgIaahhxIw/XUFi4wAqTtJvcc+9LkdYKTlWpJX
zLroGFZ9FSwPJdqSVGK85TAsnqbKM7aIzFxskdcJVXKVYGjKIxr6UHpWN00iU7G0LxetbY2M8qjA
YReZls44jdO+xxVOGxzdBQQ3X+KT5BSz9h9dys/xwJnHxczf7SQuXj1/Jj/4nM9bAkW731Db6sKy
dpL5ATc/CJ3Zq6bCNcR7cB/iOu04zdXg/ZWEs/GSrVVLnmmosrFwu1e4LRUF1J0J++hvTpth5sfN
5mJxstDViwIrIiMLdBo5vRlYo/5fBFVxZ3AhKYwZlFbmMnSAphrlAEQ9FQzLSmrSlG0w+56+U2J2
vY2TyXCMHuSkIXCgRRzTUPfrf9CnLHu/lVffntaG585gn6zq1hCDtrXJsIdFbasE9ZvixnE8qjlL
m7vWWF1/TF9c/QA2PR7eYbjZ81pzusX96RTe+e+wuX0UtGd1LLrk6FTD7cveYwiZKXuwg5TnNZ/p
Jx8UxDEXVSWiFo0WNKZN9nduF3SYrKTGcM9OVx9HmwJUnEihM0+jnBCbrDYdg/HIrinkhUzN92jt
VsvaulfOd0NkS+SfAdEXd13wfiB6IM9o0BDRmrMRjY6SZtkCIYN2lJkOD/LuhLw+eDqQS2a9Skhw
m/uz4jenTeJP7tZw0udw+Y6IZvG2xkoIS/LUBDc1A7NSmrsDG2mrwcUAfBsj08WTqn2Boa1Cgfvl
TV48zcINcx2ZPJkkesrkEHxe2/0usKdoZBJiPMhwSNTxea+sbqQ0/9g/olneaA0+UZFt/f2S9QnV
Lx9pibtYiQxkUSJ6cvQ1vdAmFHmFnUElm4ThQuqScpAyunH7Ya0WJsOn/c9UTVSvrYevKye1xhPA
64XLQWzDN9tEIKA/yUi60q9eIZjmGUCGsR6/NOHkuPf9JzGibVaip1pJe+EoZbAg6k6xOw1vkFXa
/TzuSgPwV2ZAUSIrhl+Xg1IfLYcOOPPCvMwosKYYy9iTdr0zMitVU/f0YZOj45pqElSVIPQNGM6N
LaTzTebgfDuXke2Ugc0T1+eWuzQGypphfRtJNJmLt1yYfwJK9+710ohAYmIHDnGTqBtrZl+00OXU
2aZkZ/rRIbKMhHspBPHHtJDZGhhvnWaY5aG6ACmuBWD+0mRj7A+5HCMcQyJJz0QQwhGWz5gj9VgG
opLVt9pxJEgK/85hV7CUbjUQqMTXfVp8ndutHaHQ6hJDRGiMxOmZeLiJSaMeVnoR1WdX8sXhV700
CZK04xy9e8Ia5B0heNygdqPLH+5adt4OnF98Dz1vZjqtGpZGUO3E3AadKxnWMgA4W4nMNectp5T3
h/JsTK5IXFRPzO0RzHWddzTKrQDpe35cYe6FS3oWBh8wgjdC1pyypeNSUUetYvIDlxGFWiGCHyQw
wwjD0VtHWtMK0mOGubeZKqWZ3Asb2HDEN0r2KW5MdBrfuPoX8t2fcGPfq1NqMQKSnOXeDtZIqLR2
17xcwJwTjnjRBDUkuQWugyfwOjHW4DEHt3caCtvMHqqKAYAvKNnN1qCRd1M5rzAJ+hhWRzkGi77V
7NC8DaqsCufaMtEa0uKiS+UBL8336TUA5oI7PMvqLxn9RgpKd9GoO0upud3ILBEF4oSHiu4Jj3cs
3RM03lyQQJBNX8OQPGNrnOkNtXV5IDiXNeX9ej0HKg3sUfxBI0dzjTzdBlX7Mc467Yotc5NvN2Sy
ehj6eINkNBVFCBpAFoT1vWMHpKSWfYa8mG5/NLdaekJKZl8+ggSlgFBUu+RIMFOIR3HDjGtCZNOl
35oF8mXaSzzp0UTxZjU3+7mOWncmiWpb7g9hxOSXTU71eeLxL1zpypZdfX9TW62sJ1r0Nd2p8/Ly
MViopKJwcrTlPUdUEZ/dev7OdC5/P0g5YaeGuaUEneicFnEUnEqvJVmhVP0hbt7DNzDh60edCJGa
Ctht0MDfb+uZPdUGMYoMWf73gnpgzyuM7BfowWt7Lnczhevh5ABgEULsVZufMBzxejJ3ExuqRvoL
YnRg3X+568/tqqjKQP5cB5hh5pn0+xi2RD/Ywq6j0gSBZXMKpPs4FZOsoPXVoe9I1dbkabt/+HtO
hWDowTU6btx2S2ofBFiudsrnf+7w1qunD9Agpj+4SVhfIIXJkzYia9pq3NKlMil1hhkGiQ0Q6EZB
I9nOOwyERLNk4R1/ohPFzUIYXJGIivL+HyzxJ3HcylwgJ7KVpD+lEsVUSmpnyY5YEWXR8p66yOcO
peFOQflQvUzP8zgso8BDa3ODJE37mdAKeRjYlTu1IXhVrsus+UVT9N0zfsNJpfuuGH6jtkkxCKFN
fQvUXNiHjV52LtPnYL4V0lMilKNlGHyRZppuR6pwzRk2Yya6BYWIH8RdHv3WM59KkGffudCnywkR
pL54E00ty1bOhXVlVURAB1oDniad9Y0D6az3Vk9QW0PAVL+gp5y6YLWh9jOGLubWvnPBq0bRlyny
SJfXYxXv+V2G3bZn/Ir4VfuBq7/pS0ZUMuS1l4rnHWTkzwo45UCbl2RIbdqztruaEkwbV7dv4+ce
Xm6eoLqbVvaVd/hiJIvCJxtBSy17/BN2YwKW3ErXlqYnjWhNWyz5LEKR1XznJ1EGJVKh9qmb+HpG
LvlcAl20O83RNcL0ZKKwdYOsPOY5e9GRn8e9mi4/Nd3Vjpstvs2KuJtidZkIgiws3w5Dtv8HeUU5
vchkgnvRriHU0pT1a7tGPLvfyflxlDFYhLZqIKFDbNmnuxoT2tLa/TwFsho1Z00HUkb1/bGMb8pW
DaFmpA8yiiJ2wXRwHN/hnqduBwVbff/YuCXMHLU+f/DjVqty9pALeGDbooVnbHPhnQykOaMzsM5P
df8Get0GyxquglfojbiSMvmMeLhd82RKPvFGifioK/dZxHF+RN50m0Ipw9LBI4d1uD/MV3nv+mdQ
gqMS/paHpuRMjwXuoN6xmIaEXruOdj78+Ej66Ux1nqp3ReiD2lJBnw+H84lMjVS3TS4lo/nhix1/
DKFBg/nmOpDxIH5HIbOOgOl4CpduV1RYCCkrXxOzpP2qFkbe9DTW2HFHKUeDVzo5vesk1FBBPAGr
YjOtJfSdk0CvA0XIRv06lIi6ydaWTtfcfVLgP5YWGdzMnXP9Xx9CUWQ96DUtI8PS+A4VTtducxwP
LHYqUjiYgTdDfDy0NTFPKq+QMcuXNOiub6FqFOpEI2GQyeME/ArjfkIkBlckqHdo6EBOklX72WsN
lL/VcrNS8oBv2h4Vt0wpc9iTbZxVl3oWFWXcQGCKcM+5nlsJRgHlFEtaINGWzqrGvQ4gpsz+fCH3
MG8ZWcytmKp7S3jtelWrqiXfONcqQ6UWGgAkgz6Q3NXr/ytWGY1VjaUUezSgwLCsqIBZbyyU9Lqh
bnuqXYsEzQbNhOamXPOCeqrjwo8zD+2DzMAFfYRstTQ8aQK5PVC0wD8yr9nyoGuiWHG4Q2Pemg6d
wsvxq7PUDWHP88+9XaGY+Azdrfj4BL9cz5uU0dEHI8+SX47caWuiKoxTWudjWseiTT7YR55cRiRy
Y6W7L89la6BmaGNUSTRExBj8NR2SrY8OrXY5prp7w8D4o0F/NoWPxIx6+6EVyNuNIhXHaAGkcxlT
cAUr+vJQCbg5oB7EWVP7xLC3W47GZQTv0zvOJm31ZRUCfnuqW3BeQ4vigF7Ney5dNcxjQk+zmz6T
kT/pcH6t27gimfZvRvKb1/ir/5zfJSFfje/0bj1nBy+XTpFB1qZO/4JwOpIXcyyzUSvrV4rOnCKo
+nuA/FMLraaZFFBsLCE5KGaJE1YQnubXXfrujPK1UvJTOXYXVdFIq+hEq4BvvgOrpNU/gkyVLJ+V
LEqiLThC1dmaUobjz8lVLgzBFbQd+jYVvyjndcgqbftKrTMpq2NOYl7t6U7xhhtEUlrNIglPbgvJ
52Ot3aa68rsetzV3rPZhaHpZf/YGMFMNxt6a0iaTeCOxiCYfX+RIMVoLpqdHffMD9sdvDkhdHG/m
XA59sLQ1r5GqGNg6eRpFdzbslL/IVkH8xmdou8YIZzH5ZUAbQ0Az+02JKeZUjUPGoqkwz1a4BSHr
WoDAvNqZmuX1LbnMumxK/8WoEXLgy2YIjK0dvQP2roKX3D3bmrnxMe2cnyQrNhdc9tgii0Vult8w
05xk8+BsZ3NGGa1TChbJkRZDbEwmlRlglFCa0hAH0XXOIndQb4cn+5hQ15bjkJOtCQ58pL1UPliq
oOPaMmJdFomuwuFu+PSsH30+bjJEvwrit6HcfzGxa0gWu4M362ItUhw6sEBHJ6aKKVyZMuzfsYj4
EvkW+wO0bkRPJNQZK71sn1oNr+4XIs9KCHRTRpxxQ/vZuKmSZsyKqSC1sYVI8JZBddE92nu+AyM8
TKIyOrFNlV6DfMYZ2HY3zqQqAqorwT+rgrUgs0wgis4puOlmmAiqweX+d2mVCu0+V3wzlGjnR/rO
ViNeOicPD3n2lopACo0flMnJaTFZlpHYCv4SGLToTfIvcb8g8m/hZzvenIxaR1ZwNYUdb8OUEvFZ
Np029E8jluXhT1jWkD04UJwPBGVNFA9n10m37hqJlDQxIuqcg7nM4zj32CmVVNo+5TI5RnBPuxK1
HbyKSR6aKib2lEGVCbolqZ8Moorgfj6LIzXRJM3a70jaixxKOTScR4xCF2IAD4Xewpz39Nt5pDZX
OJRj35x2JX9puiaPbrE0oayG+K89U0adLRdHUqrhwYgOmw7//c2Il4txLS4wp4g5qaH57nwWRYc7
m+MF09+ZkHMWoGXCmul/WbyxvEyiVb9Lq4OaN2JH0qZwUp3kYV5q4ilICmBteWGP8ER/7XWgKuB4
PsBn9lOVFSkO3JJb0+yIdFe42R0b78LggCG5sW3wXbTn1JP2PHUNaei8q5Z83s65WwvzZWQvVp1T
bASuNSaOm6waIiE0/aVGNnbjMLjeDbQaYVpWQ3cPGtDOmW4QcADjihQJq8QqG9/3nh2hKftv8Znl
QN3spMeiFQYwTEztvlAJ3r3s3fiqufNbyqDz3iBJoBHFBxIRtnmSvpyMQMtqXZuA0QkX8UD0wnHA
KWdXWG2DSk4VmSmDSft6V7fCWsiIOEJJFoO+V59G9Lu2k1Dg+Zk+e366XHMAHa1VErUHAWii+xZH
Y/nawJzeWuJtOxOD53B7iyz/6gBPL89rNQGnt25eNZG/Qy59qiYRQUrfjXf12dm+owDWiTk/8NKr
XH7AolOayMwGf/5OAXcY4L47MsKl5TdSz56BLZd0wHGe+3NMD3lyA/puOzi/AFa1Ycq5vE6krw0V
jr+Rmv1UK8UN9UbWtcDHq4voi7rYmYZ7Uf0YUCrMh/FifeWK+YuyUfn2xqF5vzAo4DnWYZncTt9o
klj2aaJ2n19zxFGpgf48IxJBzKfvL6AR7ifdT21+SjI39KmoNJjNWtNa8Lthcmfy466vu0XBzlmm
oW0w83ROIRgNZhxTsjgCxqsCt80q61MyuicsbmogQhTKPW1xI5XX/WnzNHVh+TWrvk/w64nHfe2a
z6BUD8OT31B9Z0be33UH/HD7AXE4IUFiKb80Ve1UjrnXRNJB2iMP+p0AelQitSkbLiKUs5veVuDd
tp0UX5cRyPLGG6Q/Q9WzxvIk+0eyfWf7xMgptrPe9WLtlYak0lo7H5f0yE64p0DBT1DBvsSy6ztK
WO7hIWmPK0RxUUzf/RvXP7QDC0aVBlz8F0gb9B+JVrrRMTFCycJHPSvLrmHTrpEWSGEi0s9WsbOZ
/dBiWn02vv4ApIqSS/Z4E7M33j0d6jvyK4/WcF04igf/qD+LYW88Y567TPkccNQYzIwhWgl+Hu5D
Xh62N8JIbynWSKggN6jB6nPDu6f/X+8c+wuYVeWZwWcbSnmLVdPKeFd5n+YN20LUExdHLLKU+8KL
PMuHQ0ARaVHN5JIGuZreWGZbeafDHZBGzRO4JDTQrILCQ3UiGlV4S6B7ZRvU46q9X4vPHBLNgrJT
MfIh39nL8/bw4C+G4hvAx05UYW2UlSpOdCui3CUkkSjWeNxOBwUEWJ4Edhbsw5C/vUwUOmdmSgKE
loeqoqb9R0ocjueUu2VJOmeyCgC0WkPIPIjY9pignWdrf+Elz8o6RGqegE1/sfnM0FVGZybwezvj
uYhL3fg6epTMvsECApd8+/YTi2cRO24i1jwDWBjkeJrdoFjJuZ337B5/YIFxVYUqneVtvWP1XD9y
oRsE+MUCB29VRFDRkvKrRpnZAzXdZZMzhFR62ZcTBmNQtk65H1+4/G9oaJtggHIEfTJTdSgpAQEE
jBP7sl8+eMVc4D45UmS5E9D8Sem0iSzmHYP65/U8ySRdpwklniHUj3N8HdAJpFhwC7zoawszbpE+
kmYnPFinlYDomRdpxEGfO1gA7tRG+FzKb2uSlS00mnfm97EhOc3KAipVD1UIj+JK05dDgM0yVzHF
QeIWlFzuTgwKavIKm/2mH0o+ZLRQrtbxxtMgW9KDXkbe4UfJ0begpVMUI55uKychrZrPsRWqNXet
iovrgVnPVBlyp0r2zQtNvqOH1ZUFgn9J1hxQ1JW1i7CiLmKz2ZVWIr6hd5h9IAp3QNdgtq7T/8fw
4WTVWkxM+NuuxOyByzD1bEd4Kx1/WS90WKIkDlMlXWgPpeRsryWYbd3C56saE8Oax1zJqae1vzOk
drtSY/+NFTjuGEYvfZli0iLN+y7fhmC68lgnV6YbX62ezc2Mrcy8A2Jbq+z4OLTk/XIYoq8MSyQc
QcY62iEqTXhGUdswvP+yr3KzLo0gDqMo4TyaFC0GYm26ujte690QvxmO0+KohN3vt+TcotxIMLPe
Tskp9/nDyERO9IOPuws9j5pY3LstnmLo8xKDv1AGGmOC7mSnswf2F/dtYFI1BFYlf0j9z83sHeDF
p/n1LScY0fec80CzD/KCyxMIvoeL7vpVK/Uj5oBUzdxxBhZF4wiF+JbSlnjoc/g03iazLSDuC2BB
vNVHJkmvZv+nd1Zt8K1VmHXHG5oTjJmiOhUqLsV/pwuKXST0M9DBNvBefy6x+obgP8th6dHMsExW
MaO9jeLsMkqnO5EiH2uZpUWqQSoLAPKQikwntrBzUvZOfFakPGmZCVl2+R73QfDgnPT+8mag/vr0
aggq56JkuVezbmcNqK84hitYGrB+7CFKyv3CnSSLwvhqxIu2K/QEaqD+2Qv44Mwwj5dZxUPuEVZj
R9AeZMqOsk7rdN/zAtn78YQ25iEmZ1Kx0UuziObqeJQttSgw8LqqgVqd7jdzpc9Vx+CvVqaXuUsD
tMmTRdfsA1j4e9533/oyNp6CR3b6S6KDRTMjAg/vu8QSsy/gz2dI6xXbF+w9D8nLqRy12tR1JSd9
mfLm727Da/bK5gZRXPZOg0xXI2gAw9YowJUr3x+mXZg5rCjX9+sipDRMKdMfFwqnavCt415K4G3g
zuXUQHxy1IlNVmw2kRgRqr9Df09OYCnZMEllKPPKQL4rjYkBf2/WtHwrNGFDzXZyHXPwI/J+hExy
yFwqUiNeJNN0v7idxr1AKE7kzux4xBqyRjUtNd2uzi4L7cpQbpks4dacX2On1NUfSX7oIWFiJAPt
Bj5qTzsgdH3FNmJpKAiTnXAr53cSHOfuC5vZeJat+/cZ21zLp40Q/vUZVaJhiOevbEtKq7e0zXLu
CcwKxju/dBURZovHEDvuOJuxtT4yajyB3VZ0CDHQEfR3xtELNXeW0R/vxkb+vOKVFHsbFwthhr2R
YVtj6qVuVkfPS/3/t1+pz24l8AMA2MTEWfksftidF4J42C3FRR6yXPjf/Cs2zVjPJD2z0B4edWwh
CxUu2F3Q3R7EdKFl/pEYw9w1tHtnMdDKYbzKaeG1EIF2k+BZvnLR8hd1WKottVhUabCj946tBU1o
PI+1ybzR/lIca01dd+GgBtYI6IPIqS8qVCpayDyoDcjl6ZdoSREGA/kDFGfjYd3kIwF34S+4SqYe
e4a4+TteOkNPDt+Vsqh8kSnsMfNXkKHp/N00J6p/FQeaAtIvMHn/AUPTRruzD6CH0Vm+QBPZsW9f
oulKmY0RfhzYQ9l0JuwJ3ObgNyZkAjpCBNLiYhQx/HKUBYbsdIyj2ShFaHOZrG0NVMbfYkgVBGcu
w92yAf2TVE4+28GWur3FdqYiZf8m5cYdxrwYQmWe1D5sonCEQu2V6QG5P29jLwlj9ccWRzm+9ElG
+k5W+2je9L6zdmt+rnnMX29pnL2OAtaBtuWVoi4UGVQvhxqr3ET3iiVs1QpiAUc2vSSZlIERyk3m
mcuaqdGLt6f1KoR/00iUCGLUmagoTdygP2lXbTQB6qYxT02ERbqi/+btabT9O2ijM+DnTv7ZbRJI
vex5BJT67p/Kou/eIcHIqpUjMvF0Tu64YOnSd7+gHS20MUUjydVaXv+g/9PN+MQSnlzQr6ZZHRtB
rNnqOHQWnLNC8yP3N57kY1AEiuNPKGECae+CSWolMYxgZ+oAD8E1HmGi5v/Wspl94wcwYGtRlMQY
bvO+UT9vTupLeEMFNrzjBZb9636eAwsTmn8cf3ZrTa/iquyN6Ft55esoecRT7UC1FUSxLWh03dJg
TDjG7g0NYVFBz8LBlkVNEEqP32o24PCkEIlYY29vDRyuM0S75KVzr91TREvbsupy5C+i7Vf38fre
KF+J4mjbp3KncsHq/edbXO0zIJ36vB4GDCYBsIakpif9lsvQCbvtrWCFaIX6SMYvkmMH2c5Ug8vm
ZQzQwoLYAofidXJdBp6/sTXJrwc5vr9D6cEs46I4myc+dVtqcMTZ+kXmD76X7cJEZOzkBL4MeYMQ
WDaCDGijj/bzvTv9zTCrbYZkXtrCkWySGIfD7EwccmKOd5yic3fnIrqpHMXKSurZ4pCE/1xDPUep
zM9+dsjL3E2ui+LWGQ2O86S73EMSHAH2bBtsAWgutCZHBnO58S+lclLfwy0Oz+TvRVkq2tzwy7jy
byFPUjKf7LqRdXjlFJsp0C7hmTe+sXqWBCUHJXZIk0F/dDDWr8Z4m8cQkprkbwe4n8/oATDF5r7F
9sBlRQSnHOTLD9hjQi4TjvvJ5TP1javlN+TMeDksy1DBVTeDQMowDydiDp7ghCcVgN+hHRGY1n82
qbenkW8ZbXxU+wzb8nR9/7z3Uii04Kre8yYmyAOf1jdNBD72ncRUBgdxjsN/fOYtXzZgeKxziBWL
frHJ1ewts0JMKDAqtKfwGq+RxLdC18p+lEbzOlMfrBFXUZC03kR4BhmuO1Am7IhxAQ4kocEXF5lp
GzeWPP6Qk4ocAIWEY7u1QskIVzx/sj6w0tgOptSpczPAHbOyUDdy24FhYnpR25hVfm422TWYnnIB
/msf4urKVANtAEBWuPVUJw5o73fHieHp9xQx1+wBen7d3N1baUbhGxpb9qyYKRziTVZPvsbv2zC9
3/7m/IxdLeJBKjneaEXKAeDnDUyliLdR10/x3EPLmcy7s9ky60fQglH1N6TbjdNZfgG/XtR9bkOT
jXF8p4DiZT2w5KPDjdNsk22fbnLEXeS87kWxWw8EpOCyNaw6EtzWh2m218NwTOCgzJdToaTRRCEs
Rdjc6E2aVVpkviUmLBGPPhrvinUpv39pkovHJmFwVHkaNCGLI3hUpXTKM+MYix0mVN5MPChJRoGI
ECO/AZ5aHUi3pUv5xEDLy+QBrNhPYAPTFPGgMdvP74X1kfz8HAdfAsYTx4JZEGGmkDoTOFdgeTbI
3PMkaCWZjT7zgfHSH58LnO/2kTxsaCFzaF0xp0yFjv/CzASrQRoBpERTTe/v0xVSsJVBANvyp85j
foHeP4tg2dH71goZneZVUwqQhKANRrZCgie8kFhQA8BYIPqDUaI7eBebMOUdkvvqTZdArT0Ys6GH
TzgFdqmWrP9JhowVRKlv2RhtWcmUj+Nz3A73QPigIoj3LWz2vuaPZLvmmJI2F63rLKkbrfB9Ev1j
E3T/V9LOIUfFPkAEmU/tdKSF5G8Hb7ybCd9axt090gEKi0krkPiFTasnb3M3BA9esy0cZY1LGLJU
XenSW07JeQPC0WvuB/Mj99I3FedhGSVLdn6xL99NivxT1EBbZ4Fa0elPugy74DILVAPqHF20HEll
pCgaTnorzUKVymsRxmesACzELPaCbSPExPQQ+rUBAqROxaD9q5J1VDOv/Te5fV4Nxg8BDQSKc3hk
VcSn17o+2y7Mb7TKsd+S0sJLT81jkoegtMYumfXpvEWl+pcSUqHYDSsbw0383iAA5zxhxnHlmPKC
lqMrdkhNaupX3OrGJflup3Bmf28sXHrsszLAtWbPRCm+5uJFjpN8QAfdMpBDy9F07xDRC8GpQ9a5
Ykla7FbhY1Fpdl6G79jIfbTAE4BwKGvl8Wu4lQ9/46BgljJ1NG/uH7PrCoUdMpxWpkgJ+qOVGgbp
F4LCuJLppbzzq760fQixCXie1YiJecr6961JwLxFbQtMyIAIyRa2R7cbAzSBODMg+ALEyipuCBFy
ymRh95i/0NpdjAagtH73Q9VsmEM9Pd/xKgQ2JrARN4wDiz2EjLQBP6JZd+lwdLvIzr8DgHI9BprM
t/6MufhokmvPJa95dTLvONWt5SM5t9FED5pjKqOCxT1KDHrKRxPIdp0yK/badgYOfOaVmzVWshLc
kTeBpOuKl1TF/WC30a/nybKOJoVm3cJ4kQTzOcDtezA8Id/woSZ8GmRnMU1Y9X//xqc7Anq4sFTx
2ApaY2vsHfYUxlLYkAS42o/OjPHTcHCk2DCxumJClwg85pqwzngZUcnSVbvmzdHr8dZkNZzjk3Hp
y95ygUPiyUCI7aNQa77tgCW6PJHn2aM7CYliJxp88D9VGFGhBUixsnQ4Hw/FIniU/lzQHDCz2nXH
e26qMbJ9IsgranaBXik+AVY5f4zsBF/OzxzVQPx3IKcaHSRQ5hxxhQzS96GDy2/HmYJyM84JfWUg
K8Aofs4pHsWjWhnfANnxUspe9PHh2QislfDK2ZsxyGj8hhqEP3CNo4ej0IBy5X4cPBB5G0hYBn5y
LUDEK39Sfj3EJ+cTsfkfGwV7Ut1VtP4Hfl30mwP6/mkJZqs26pT5Ava0Mh6vy0aJpiiu00yMNnLK
P5fbroixQipKSVP358TuNlckbNVD2erFZ6fmA8UtaHtW/ImzQb2zdqg/tzwwafweNS4jh8cErc7z
FkSzErRy2BPgIH0mbgKtN7Qq10MnNSjM6M9/EYz/oryD3LgM2CxOFF8OFTKBwgBi35FcD8UjQKgh
SFOOM5mSfHqb26Vq9aM3A1d/yPKd9Z0oFZO7XkzgCI9TnnNd5JieW7+3mtnV7/P+uz5JUq9A69Sg
d0XCTfSCiyzl4K0HMcmHxeWDJorspR1JKmtjrMwfzoOH0veHNJiXVg341QL3AoyfCI5UoSLPI3sd
gmWoL1/nETvutVfNTnZ+6pXKyc43bRnbN51r9++FO6fYNHORhEQ/R/QqGgqD6MFmjl5Ruq5ZR2o4
TihFwUTCHZunfjuTjJ27AkRW5t12Z2msKjlLp0xz4O6zvciU0PB/AeIAl5hVmZTy0Sn+IqtWvGql
IAIKvtYBEp98bzJgTfYDhzX8SYgVPPcKRPxBDn0QTBdQWPbYQnkbxTRUvlbqXFQlsZKzGDrdQgDg
46RKrEUFBgRMkmEg8HGy9CHI+xWcNVya8t+HIqYWUOIWqR6tofNwjWRhloum4sjBhBtSSJvVuCXj
10DnNGJkrnO/OtIk5x/yGh4b+RNP2fLmWgTWx6V8QfkG5S5OU77DV727/mC9HO7EyDp/Rryx+xzG
BfbdDowb6H9zv/KFklSmLdaDdxtFxRDRqD6PKArrd6ae9k7jKwHENqkvkKzhhpuYfas5QFmCm+JH
cHaH7XIliWEc12eQqkSlwUNxzsTq6uBNchdZO7a6Gt86yMuoFBijH/EcfmXw5ngcN3zHGRC8j8mH
s8x6uktquC7EbBAMxD0Gge0iDh7axgIMEeWnS/yWuW3MB5BUPFUFEZhSnAYdCeJK+Il0B0Tx8Hfk
bNVRdODq+Hk/uM/qro0n0fKtVBVHyF0dPkhmsWYgUnsy6Eg+Z3n/zAEmsle2p+Jpe6Khbe3eZtX1
lYCYn+9X2nxdGAAFj56RYDHkaF4qllkYT6Cw77QRgB2bshTEkf58VCntnnWJswNS/5WHlLY80+jZ
DFU6bgIS1FaUKkdrvMNKHBmvC8FURSeS63UpqBz8boMrNMk3tdm3y2wvZB/naLueC5LzSiWMFeU9
IG7IKP3V6v5ksECVQIWJe37e4BXe9rZQXkN1fXLyZhZQUVwJg/DWLhVvPtPb6QpKMTgyk9OJj/iL
6/EDS+xN+rpZOgaA1zm7tl145lqopFAP2INpIeMPG2sIwk0alBlYJjKiDBwUJiRhCFHRSAOgXjH1
BIOr9GcqujF1/Eb9fAayoLkF4c+oNybkYt5kOnxHDzpo/MRXg6cRjc/EybB6kZQb6wXoB/NKFO0x
xBSO4NTG2mzbG6xqPZwdb8odCDHkaI9g3GFTJA7uzsng0oyOEvbNSB7Njj3dk1zIqSTGiao7WK3R
EHR1NJnnL8CPNukbFeqXoDHZkjRgFpOElMUj8YOMj8GulkTKKy+Tf3a3GT8ocNA63Mb7CrP7UGuc
leivSEWjt8D3rRUjkFhlkzqJWjf85m4CiQxpBv9KWx98bhi1KHsRy4pcg2DVxnIvmW8Fbhw5q8Fo
E6YknFAAd5PNmKK8u1p4S0V1cEd1WYOxOPklBb97Gk1uPrgln15ryWgMs/XWRvIwji61F1Eco/NM
4at0prM/IkhEgeogn3/EuL4SqUYZWmmAKEWh3av9djag8ufQXWhsY1iOtx/NeUQ8DgQXEV3EycfM
SpRZO03bUIecwYgkndhZtin4O74RavaszI4VyQoWPOBjEdWTJTsuuywkHfe249Ebl9RNFVrheX7B
zlsphadcoLglWRMNynG5GvEiYkc5MA7A4CG0asLsZtYLHHTJzb9QoajJYYqKAQ6NdwjXo5nKaAxZ
z7KnsHfJzGr5LgckYbOCejPnUsndoTIYoIAAUZxcC4aKhh+VtrDlt5R3Hlwk5Up6LWms74GlZc5K
uA+YidvrL/2XYMbdnCgoOXc6MQzls/kxmne0TynID4dfKYeyRsp1+krdRJ2BK+gbo3HTpPk6bTXl
2GJYQI2OHX7K9DwHcBvISKqavDjCQhNhd9EtGCLPCPYB8YorPJgzMT5NvpjpKiRJKhAEl9oYRYZb
kYgw70eKWpAysRGUFW+yx8kvr1jrcGGH57vImYYWULYuLr1KcAF1w2qK9oA+kfZrh8VBuQMoU9gs
RKeDiVbNmssBWZhMEtmuRJdTtldu7cUgqio0PNaJ57RENrEhhevy3ccqIwxeYYhfBc7sqQ2ThrVj
yM2uTYmlRxV/+owlA2uts+MiTjtY0JyP8hAtLHMSKCtAGLRrDIwIFZwdqaPz/AwDO/PW9lCbomn4
m/GGmMCLCjyB2QPnAEOfYAoWhCBwpyzjNlRKRaNzuZrGxdIxIBwvp48Fc2DJdaAhSrS6v95FlmOX
ogRvG/lJMHWPJkrq8JS0YiN2y7xWk2QQpriEBulefz7aIidnF8Z5qTycPJznYnoEESAqO2jy82sv
8S7UkKe1jPk+A2b+5dy/ZAW0UXIeIUDy3AmG5/GVfjmxSl7TZhXjbQFCRUbuaAEKIOSqFYaFkktI
7qs90uyoCLpQiVIZn1vFZfNDhg0JDgdghlkByvCBj+ZCYL1pQNzg/07PO297QvNF0TRlhaBFf7fL
AKtbHX/wVkJ+JRDbKSxYh1dyefOIi+5LhB7QBgOh6t9VKtdRIB/+idqlRif7ffpFzWN9y1eCzT+h
a5lCw0oGvhLQArc7o9iB/F6xe1ypNeOmkDzkDF7HDZuhsPcGe0IPcYPmPTqe5CEBWkhU97q022jd
SxalSeRPw0mHC0N+Ti6IW8reuP1Seb9y/K4Tn5fuFDWs6DoreF+SeYeFwGuCIBX9EcZn+2OGvHy1
k5Rr9wXDwFGz2dpJWdbWtSR26OAhuTfqPtHXtqy1q0DNTNFPa4krvftSG3MwvpaSOWuvs45Z1Thi
fOIv1SmWhAaWcdaQNVkvRBKiPtt/YjxjE4kLDzsL8UdkgsQi2TWPnXEmnC9NZ25Mzrf/LERnK/gB
vb+KRThgP+ZvdpHUg6XhpzENTfI34kVyIeOvyx0Ye/WRG49vhsFz3ZWYsWXUvWlo21mqmhc436Rl
WIBUwIWNK0/RiU1Ezvkdspv798zMAJ6UzGhwv1nHswNMRyJRTWXiLEfxKuFfLP9MdjYLjpusVSe7
Ld02urN7ozPsc+fG/ugH543NFIqIdwPPuccroR3CB/aZype3ZtptU/EAj4Zk0YqPMVY/VrGGazeX
HjBL+KBVvCiisqhk18SLzbhjo+2TAYiItWM8GOSYNf4GC+IMk79XuDbOPBvhb7tBG81uX3tc8325
XHtXE9iK7WcjvDIayokwZJLgeGmisUpVjrJ5s2AjzEt/D0060OdB8eTCCL1qBRKGI6h82P8IcKS3
W/cY7k/x/DhYeAoHq12rMTO0+2RJzOfqQTsPq+f4Fp2yQSvC1ez/MkibB4bBricusk4WoMVCxTmx
sE+6PeQo2UBvHLWW4ZyB2E2+l72ano1PnbG5P7+y5CNw329CTlTBOHKZH+qrJq4F7RX1lOHG9NbL
ys8uiLRfcr8VqclMP72KQFDqjPP62Ru9G9ePpY8i8CfzHImyWp3gjdM+x7hZvq1rwDgzcmNKjyXc
3WuWLch372sWfaTl5f4pyAd5D0qxddQ70dWoBg3Dvc4/rFgz5B03YtYtKneTCd1frjpBeP1RHidG
LvuiD1EMeFDfYHJS99906dMeOLzkSreVOB25vYQN7wJ6yBGJ2P229xUtqonSaAXuxWsNEWf7ctYr
kgYSEJjV4Tsxq/ChiS2zUxMFzIHzCgSEM+MSsZQYvLrUucTtSGbJecalvK+6woOscY4h+LuYp9h+
kbZTG2Sqp6I4OBtPhGnpp7VVr2HL0xhE4xWQIuW+H1XcsGP3Yo7NXRGzrrvCL08uYDNfutYwXTMi
7ElBVsVww6Bv8GjJ1aMgpEOUJcvCDSPchFc3PXG9aFmzGJ3C89CE6wyKyveRBx1sXkLplNUNa8iM
ZBZlkQVVZX4oR35sxLUARxXjTwLkJwt6BmqyzOasTdNHPE8lZUhxNx1q0kuVvec2P3hGFHddEw3W
IHAmizvY1f8n8ae2L8KzT1pu244IGVQ3rX35sErrs58ks8P34CTGtWiJ60tIm7/1TpgMZ8MyfDhr
+8RUzSLMTJGUPkzS9T/2RTMfPLEHM3LaqcrdUhMmwIfLsOuqSu8ROpc7M3HI8AEUgncAf42WyOCu
eX8szJz0JBizgMnqExg+xJTnFWfeE8KsJpV9wvzRwVxa5yHHAP+NMgnKVyYhaM1LsuWGUFlODET+
V2gSzo1CfFFAQanQLvv4WQGQ4ZPN5kTr0F9BZMBPghlKm9yvbBKWGy3GgY+yvLyik1ryOizwl1jt
jiNFvuY33Mp1bJpgxX9IfHP8qs1n5Z2tLO8Rrnf4shKTrbNsOtZ7jxh01nr0sLPaHsUdWdBg/N9Q
1cuhTWcaKDlTZu+aUumqebnhZctDp+w4BsPNTUhAorVTM3P2An/DErwZn7wWOBMEoihM0WgZIn4n
mKd0U9bTXurFXBjTpYaI96ijgO0jZbgfAhuWzOrVJNgZubAWXFiahye+AJiZOSgHC7x9chV5UMf9
5lvq7vflSBSQM36fp81qiZQ97YG0q/3QzbbOL5IdRwdhffscmDuk5tmzR++dAQGOYUJfd70wt1eZ
gtUrHwS6SIX3zgXLXyNXT9QGcCqyE4xmG6v4l2BDp6/NsumZBwgzbsQ/pgY5Roc0CGtgk1Ek3734
fu1MBqW8Ld9XBxfWA4pmQKkzzj+Q1r1QNk03nMN/6ZX3HcTvenrvNFIdVIk6S6F04HSrVzszxqB4
GU4pb3TZgruJTb5rToRgniBvhP9lFUs+n/0DTvFsvKps7i/QHAq/Xp36//0sj2RLa1LgF0Nu4GgQ
/GACZWV71qqlq1fioQyWeBd9xY0bqv6R3DJeaIeVYLQ3rQmYyScd/XO/G8ZjUhBrN7RC0oOz6fvA
fXV9G3J4p1MdqHAetTWzb6f3Z4e7yX45SNf4hiaemMy0+Jrg5kNMlRhuBJ+GT7LJm4BTXGT/w3Cp
mPurskSnbbaBpJ+GfJo7+ZBkmdUYNr6SkqKFOd0xzlteRoDtupOeSXiOkKwPIVyl5KF1rcP4HYOQ
nqFasF/mbro7xynVyKNxmFKTOwIOs5e2dR9eD2evvM6hbQ5bSIiyFa33DasfhuS/8X51WXz9pL+d
hQlw5YYHiQOmoU1fDU3oDqESC5mEAJ9VtiPLbXqF0EvGO51TfIteG5q2MU3PG4mXbNIOYgR4u0iK
FCWOm0GsiDiTAvOqa3fw0bfSnOPn9U13WCKq/57IJ+pIWl2tEgGfJbJYlMZZcRjATG42Ps572Aad
R3oKTcDo3D7CLxHpi3oEgYxQcWnobq9y0qGr/nX76y726pH6MsHKiHHNPRZHI7+MCU+OwctjN28b
e5Py7hQ1KJhTRQbqGrHk4r41Xwt3wdPlJHtosDvwwyhnl4Vujhs40LJmRznK4rWMAQKCKfKjAsiD
gFWqm9emDOgAcjF55Z+IyuOCeFC7lPKgCc6CdIS+Dl1S/KVINK/ECq4qBERKPZBynK3J2diJZynu
JleytNFohjxxh9ESTcArTszMA/3jM1jK7gw4teJPvPNceKF25y1NbCQ1iXuOxuJhyFyBZ4LhwF/h
PZOs35XqrTfCGBrd//zfTJQYg3Yr+Ml5Wrpo9XEUl5GTw7m3s8jX5LXCzakoNM8gvNsa+xwryxq7
O9ZnrrJrg10odEfmmf1Bpmk8ptZNKl4Vq+jl4AMKJEKPo0+nY+pO/MAj6JpQWx2Rj04iDkOQ7yc/
eGR9MzLluGtCLYZUHxOZWpx0xj2ImAEbC/o7RWYq//uK0A69iQueVNd/Ft6j2ArOSTKuA4tD1Qry
xnGx/rxuucTlS7D+ID4HkqiOm4rZlDyHAgoHNAHqtJv8m3vSgXM4If5gFarzfZPSijr66pdfWCq9
nh0PDZ69Psb1+tPpw576sBHTGPQ8mr+p6wvT1iZTc2uo+m1JQ8j1gM4o4Jd1kkoVvK7wIwCSeuCd
oZHsb7i6GSCnmsgLVvz7sfP4JILwinuKjOg2ctQ23KKvwqph7xc6YK7/DDOVEYZwJbJ9D+eLEIp/
CtnfdPTfe4gjvtnw1xXv99ZEwn39KbltxxKs+IgUxkwdsf656ABpgZpVINzu0pKQj5fqpdiKKv0Y
1+i6jbJNY3Zpi3d/c/0Epi/WRKgJIReEkqGgb3Sr+sIvpA1vOdQYn1/K+sVyEFdySgBcv/GAoA6B
+nf0c6ymHgZZoe7XB7ROZEhrrc8e8Yt+C3sPsF0+YVEETTIbhToSRSoSlWlU9u4FssfiJUWw1L1+
UPR4cFa7Z6bvW4bxml/4TDvfQiRlnxv+ek0vQqazNIa6JNHB9j+ALs9qatFwQHmNgxeI799G0InA
aW+y3gu1WFINWi80gmeHuqvFs08kOxtN9Jg75e214kztVhnJ5eqBepOaBT8sQHxE3cLw1S5Y0Gru
agxUmH+f+Br3UcXxblcxEhnuvsnHkx/XZvx0ZsnMhbQUy8isr1tvCHBv33rMOzAnd+8HGSVwA6jQ
kDlsVltxQwBTL3r88XX0Ucl31yAG+RDW5WA2u96NWWo5iJaXLxCVYDIkhFD8CdgByD6mo05SMFRC
C7LGbsZeZm/xHEwtKeQ+rNLl+OZxW5ptrGQBXI4zqKvYRMslPY2V+t/Kug/k4kKA1vcRd+ryeZsL
5Z9OIfUrorTuwPk9UUhPugnSZR15s6X0GmlXOctD5aC/W1jN4cDZUdV/brWwO+Waa3eBcBkvmc1x
zQ2urNKfpVDXEkuJk3VdON9Pk8+sxOniQloAocq7vCCXLr4HCfyWcxN6JMbBnfsBbQyO6XI1N4Zn
6I+LhD7SsznRQgJIQlLqgUHOn1TIOAMJ9ZDVXD+BQvGMlqLBvT4m3j25SiCcyT/a758M7wARaVN/
NFK1jDnOzKVgdVfEr4enPjAh0ZXjQSTvLKM03MPcHC4jiDR8mnlLUrKKUVj6p/6FBWYkaI+Ym3M6
ltiyoX1FVrniUiKSAoP6o3pVpcUzrK3lmQA0/d2HQS1gjq3G4BDT0GpzwNw68po+DPHoieVvFylT
Dg4PhBG8to+N2ZoKlmQClIjwFtdiNq80FFLZdOvlnXTff4htC5zY2i13gxZktCiSzPnIBlqb3XyI
HmYxDj4z3+qcwaDODgOBtx0+ZmKM7wdTlK3VQM+7BN3nxrxCDnXMraZc8fwTjzRIEPQeQSjqUCuw
o4Y3ICo+pgUQrUrF8sIsf24w8RXYzn/f5tmxqWY3VnXRKqbjuNcihY0rmdmVwJUUiTm53F5TI7/O
WqpTN4W0wmd/TCDY0yat2e12EMKzmUdk+rcvmjmF24RS0M9MGmnKas5SCG4QAiGAomnHYpFtQkHh
On8fdl/RpRTxn8/3DqqeaaZTrBsOXYCH89rUh5dzha4wWfthE8wa+UK/LB1iupF2bh7IqhhSkTyD
dDMnEmZVY7+fDtx9yQQGATjU1P2yuw2ffmOcdFVNyOy7up6Hw/KumtOGhZQFATdpUMpUlibwCFVm
1PE1/EvCxWoR2RWR6mdF6SHWAasQI3PE9zp/2ILO90rgFbvcjW7CP19ZSnyjDTb/OF2eXSdwTmXk
LMO29NMfkfnYMhXSmedujmzXrKodlPM5SRLdtE6cjXN6b/TkbtgBxxB6gSimCPW3rTgLnoSY2TpY
w3EcPYL2CUZFcAZWtMwdPlEkdWXU9XDcqvDVUR8AJrUaJY1zt3hJ0gTzeKr7PVdROF7q8oGqnWNL
fDN9FkMj9VlvhM1gZe/j+Y8H+Y9eoHNJ23CKPEGbEqNix8aRJQeH+xctLm+hPQnQppKTQRH7suJO
XaSFrl2jo1n3JCeNP7tE2nTC/OPSiiscCdXGQujyK7X6Z7XYdbtUQJ/jCBTeUflKZxJijX6b7CeB
uy+OXUh7LyNS+8Lyow2xFDWFqTKe+xQt7VYHqUmHtfnt/3TeXskMIb75ftW8PrMlOI+qyZh+X0I9
zetZ/eKmY1y2UFMHIKfA6iD5lE5IMkMg9pbq/lpkhfO5Sw9kie9nwYMJ9xo4zPyMEU4Vkb30IBZy
ucHIEDJLXutdLSjR56ckmiV25MdI1h+b+2z6dZYIp1mBkGmz6jWwNzuPWED1EcVrZKi39ZB2Zxlh
avWw+BXQOz2LPUw8PUm1iQJD02uGaG9UlwAYirn22UHwF+fmgtU/GDJHChdHqPuvIGcWfP6afD9k
29ByNONqjgKWdNWU/AkElhPHmzgwACSM7pY2QwF6XTR107zTcpbOoBhCo3dllGs2+l2fldUTHG73
g5HZZSLerzfuqM+3XOppxVBn/qbiOm7ebQH1VDq4ldG75bMx5v8zC2iswSgzpnNfxlKKbBGTv/6o
iEuEl2LjZ/DNt+WcX4I5z3iwtr04Y5fjwdM38LQUZieiDwKOY0wrEAbV9DvjWsr+RWVUQMPCknPt
MgwHzqQIzlDSHltOwZ2SwRwrm3v00wVA9WFKcOkuu1deQ0wjG0eK8/hD9wTkhemPg3+K1rSPWpve
0AsWVzJ01cEfYjZXO4JTzMtedmMii3oSxtzg+q62p3E6DctGQkYjpzhqD+PPhHY9T1szNRY2ml+9
UkKTjs+NoWRwc2W1t/b6qF/Swf8DxLukiIuSH6vv55yoK39hB0VDHH3GHomytUVy6FhaeBpVb7Wk
MKCxCZEd9NErBPnMrcdw/AZX1QBTBLNxyfbg5juAxEfQhTuQ5TYhADWg1nBXGQlVyx6JvME+PsiU
yU537yNMfdqe2HxLX8FGVQvBeUWLNwOYodOxmNQjqLIDC80OjdT2sAG9T2sTw+CrOZjok3orWKMn
wRb442shTgckPtyS2BLK9IXxElUJwCFX2nYBqkuajo/9sVbW4602cYgWMC5SbSJ3e+HGJ3D6FWXq
HUUZAb1u/70Pq7CDyU/gxXncKoMUYKbAoOmsP9pctc9mPGszGeiZ+DklYigeS+pFneJXTV2PO0vm
GBN/KFHLcF42T5EUuHMRX4ve10UOkFbZs2sJi73FZ9XgjPMuTtt48YwF1lLI2ob0/n23Kw7M2F0W
Up+Mr/P3bnvUX+tecSVo8VaX5bnUrBKb5cOd0D8qEKDlHkWeFHuqLHyrfcX49MIqUv4oLMS0dOi6
gHE/QuYfH1TB67iHRoPtM8WVGR6xQHN4D9bLeh3NjKiJCx/BsDdfATQmm6PXcMIwivGG7R4avQEs
eumkptqy9Qfqcbqet2ZPbaYRx9J6LR79qTc8ZgyHOJyiEw1/OEnb+ufIMZ/CzTwIPK4VY2wLWQ06
qJGI/Me840DD3hqq7zqlCZG1ByJxpRCsh3NMmYhIzEqTztZFozGX1WcIiD05iscJS7BeOzO1Pf7C
jIi1K9KZiOQZfbImxAY8bpuFvCa4QKqyONYrS0lOl0Dcw1XK1VTdZi/nWOrM5f2NrkDFbAmirBDv
y/Ky7LaNQNj1GW0ig6XcpI3WVDodIYzaeagJstlc2PbvaZLOkRFjDtP86WiM9ppPHWXb77g55zqw
e0b4b/8rchLe+ZfyiMKrwI627NCY2mek5qulr1ysxReHanzWmRArjlz3MRo5qfRjL4dZMGXm/QMI
w79YjVtbQVMLLWFkfd2qNtVLzR0XttsJap2LWj4ygMnvh+8slcQzAbPSijMhF5CEC5BwLPqtJ/Ai
1fCbtKUf7F4tOoAb8DkB9g/edpQh3LP7RV++5MZbxQChqGjIRjC26FHFENFt1Bo0L9yEHOqO5Vzz
IA+lBhFK5kKha7tUAn1EFatGwD/kzXW0fMsJrRUGTi2evglX9FIT4ozRu0a3wIdHMiaEjqsuMWPT
dMfjI7sBUW966EgvC43VooC9ZuVrTfOgGd2vobptCONwasuLOJ/DVtS05Ls8ai0mG3l3aH/QNaNj
tgr5WOyEalYujUR1zhSUszUUBB3Rczrio0vuvNcJQ1zmUMbUN1XAQa12H7gIURE+/Qhq/X5ycBHW
GoxABSJbVCoBB44iE6+WIL+TRrtK+4R7FUKwIpqHqoglMdwmi46qON/hzrHcSBEyHYSkJWQHJVcF
VgMEb5eASyY+/WxXtSnXJnLLJsCs0KcjUVcq8LsRWte9lCZOk8ZWqhbNb/d0OHGbg/0ZHn0HUj3q
WeYOzPIrrzJ4usHh3pu2uj6zdYywRDfE8eGRWFFhCdTy6AV9BxPXwVxJFeNT/X4MHx8f0IfrAKRh
1j8AZpWCaYIREAnVJ+PM6JSB6U0+luix1TXOht3k52BEgalCYWH2ddx+WYtm8EQGrChcEBcteyMg
aT1jFbEGXi4hGcBBQGQw0e3C3kTFtIMdD7Gz3fyorwzK0bnuir+hy1W7jrOsiJGby6E7dK5qXApj
49RUd9390z34DqiwBkGYRzdfBN0THjdJIHTK7SlZfXKmrkFNlKqhVYuMPnsyK4kGslmAuc7o0CD+
hvnjgmlO5K6W6QMcnYvjRbZ6/D2txquOduRdzl9Jm4KQOyrmkM0YKp7POrGKurkyWiOyeJzbRJaS
o4OGgLvIhnrDn3YwDCCqHN9e5PIivF6g5KbNAaSTJVsR+scATt9f1yJrNo7E9C9p0IAw4U2O+6xr
ECVVLHz9gtlHGJeTUbX7gW/AKnUEfBgN+rI/tU3PaasoP888s4C+f+0H5TKpf8FimT/oQ3DInHLC
FjisIdGXum8XY2zOVw15RvAaQq+3S7nW2J2gx8s89GnoSUAc5dnJgUHfPWrOgqwmTn3hgX/OYYVB
phL7mhEaGea/2jf1J5l2UW/cF7NK2/D6tG5FRfQaItiNjeSPtjBl/Gn0XzUYunaXCEQetXtGI3fD
HqcZYK8Mm5sTWgNyb0v3Kc0pN8LM8NDnaoe8OcHA9BtYUJHCwrML8HVlipygAQbAV8aUjxnEbktl
zvwIuCgAbi0XsYHP0+fCJYrBAy+wThffqOcNiFJ8d2gNq20A/pwjXkYYRkYpqmnwHXufGpgPcInZ
cuTKv/p2wACLqK4pKrjyqvxvGB43Y9TzearEa6mrKq2DzWTjpFylotQu3HgiNefrrluQjYBotOJv
noYrx3D3Ia0y32La2BDtYp1CuD323TYzffJvo6Pt2OXD1ssUUzFoKt0BYLz9gA7O0sMPtOVDztgz
T0WtyX5PRYeiPVkf7o+xWyPeEw6Uon2wNatZqjxvsRGUe0FgZQIOZLblTfWZsX+cJaRYug1C0AJ2
GNW8OVQx+BEupY76MP5KYerN5P+DFZ7edYEh/ZlPDsRFbbrky6T5/TyFnWRR3gR8x245oV1HW7sg
m8r8ny/iZ7kS8iREUL9oSTc3B+fKaNIrmI1/0D1EgsLeo2AhvBycHhZuI7EZhST6Pnqo52LcZ6Dh
kKbAypiM/L4RoNf4iLtyb47faFISEynNGiDy+fJbYtHE5mv9QUEd+DasdKU/Jmw0M6KxfbZHotIQ
Pu2BLLd9/g3iyF+L8RveDFBsPldi6824qa2K0UxKWMVdq5dIFB7hhoe8JaImQwO6wP9neuTdJXNz
pZVfmYLBngid5fbFp9tSY4CGZ4QFFJzR/mCx6KfxTs9o9Gd+dsAI8Ve5KtKXkMeDQV15LzaqGtHg
mcb3HbcZQ53g2iku1bpqFSMegXUpeAa4ld7khQSyTLdMU/W9vAlZjyEeV9aw5fotHHMed3op/Y7m
iFD5UFKsRJnIY0bHRy61QZA1iq2uvQ6uVD2TPIA4Oe8MjPmXLBkAVviIyoZnVoI6WssmWjLLeAt5
nBN1EW6fuDJA4yHYCmHeKjgWx0hQl9lkc9balO2OBEE2GZJJURmzrUy8ZoOcGY3DasuYf9FeFD5i
fXUFpjMtWHKj1GUECfobQnbyylbyT4M2T0Ee2yiYSpddyOo6apckb2+8GZLF9ubFCFDyzY824j/M
+OX99996NLycgPY/DUVS5nF6EdlfTn85zJxSznSA2YmvldvPeeYQGq7QhuSfQB+yB1arK5iRkubl
wbbXrHMK/BkC6GnloOzUoziK6sFGU32Pgedqf5cvALmAHvrzpcLIHWfdsEnrma+93IDdgm6Fud9A
voziDg05PSXMJWTkWldE8VipTivAoRKoj2YUZFuQ+VodkLNaJApy2atNqi21Nm0s5DPOetRxhq+N
wEesvzdNQ44tbx5/XLURtRfcry9kq4UwbCv63smKoT0hHFwtA9B4TdJ+K0+2hBgHn+DCskzJr3eA
ymQTbtAf7lgi736EQAdhaYJkTch35QMfc8S+MqnZ2UwNH5kPUz2vXSRCEk/y1gmlo3wkMuT8n5nx
WZdkXmYAdNSCOG9a+PsIVSbsI6WAY+/VzhZz/CHKacgIxkDZk/evP17weEP1vC9jHGOxqC6xObI4
g/7a5vk8aqtcZJ2ezWAI9DyEpB79pjCpyyEMsWdzCcQ6GMdyzRg29B9aYwZjb75LEfKboBFZi03u
igE6juntyewabowCtbnuNHskPUR/gPo+UlEJBZ782FJnsOhfGR8v9yNW1sGuSKlrkBzlDEGS1Lv6
ascXkwfv7ckyj6u9Ph8NDinCQ+imz/sH9ycy2Xg8XCJqq1bxpISI4Mptv6FG8RXWm1Vj9VnTZMdo
JnLNpwzcEuW73A8BsSFwfoP4LOylmkAjcexibQidjguCX4UM4yOlxg7HqT6dybFPIvVbWACApXWD
ZHU5Z1ExA78w/Mm4yhb3Tbu0LuzTO/Anbb832Ba7ykPS6XjDvnPJRWgFcQ1u1BNd16S38j6yZ8Y5
MJU9E+kLAkcsBTE8W/LKzpiDdut9mvf7kypdxNNkPp/UhLedjbFgkBIOQxF39MihHBZAiOrZ91GH
UYuxnaSkNvrntnSV1HxpXHORpI9hgp7jemkvzXKA/H3tQoEfY2RRghshBZx+WloggjNE1l/sy8ci
vO1P1qkA784mUSr0k761b59ekdbY75zvQZdvH1oCLmc9qf3inEQ8UuEc+rjaf6EWtnCfo2Ai5LDT
tqvd90rvMY6nVoiHrF+PUNBZSF6zGrk1A1xXVPx35WdTNiQdCR209jTpJq8/u/f15ghJuWIlqDp1
B6bo2ykGwQ0UENSr5oYrp7rjQHSDb2/8OcuGPNulZkgbAu7yw0Dh3ApmWb6ERvuVhVvDpkrp6vLG
d66ft3xa7hvKxhLlfiNdBa+CUCjYI7IrnPIo29nZDf4G3KIzh4jef+YvsAmBa66DQEmc408Rrjjz
1VZXBfg0kRWam1A69ze7a4JZToxvbIwYyTDuZpNQMeeP45UgyVzM7esgVKnXVJpD6ydPLDjBaHbr
CvAxohecCC7F/qw/mnkOqJHEMcJ3GvQ4BfI5nx3jbPfehhzTzkMTgh+dejPlZRpahtTt/ltAhgQv
8zY7UIY3y6UUXksEEg1rhazTSLFlMr+miaRTPgkABT7c8zpwhupgQ3dWaUW37YDz65MJt43Q8a3S
AS1+v8IvHvwnbEYgzbEcWXJcW/biNcgeTRnLYsA40GN4/oAahexPZdjzjB8kUsIwi2MZRD+w2Sof
UVe3k/aYkXoPimemOMGA+5W+PpdmEB5Rc3OABMHtyEedCW0s7m1+u3foPMFUft2RLYDWt9OqVapE
oRDe5mxstrmwuhOdoUDxR0CSMtJy0SHJf61TJWKHyGRyevGei5gWYjidc6NPeVJmrktuj2ErlV7U
AjZ4nQuMbrekcpfaN3BY8YgX4HMe9ivHK0eDsiFp7eIVJgIQB3/ZSvETI/QC7JRvt54e0EKiA23z
3or4RzTycaM9g33u337+2jK2OAXqSiAE95/q8CRz/xnDXGdwutOuDNeN/5vaevOxzribVXYyOW7g
vstpDXYuCy+LyGwX4Ly0C9Z9ixQD4fiv7k/2CBNXpuFixWlsjCWg8rUiUVtE6xnq/G09voEGey3B
Z6AiahA/DNR4rau886kQ1NRzkymHtCo8t4E5XKSSoV+1M2PcBXtukeDJOPzEO+bCvSQzL3If6hRf
esMj8HScOe/KvNC69Rs+uGhIwnrPOrxaUaSGAJvJEib4jBAbJ4aMz39ei4mrl0BZNfz65FWUoP8d
Cn2HyJ0nZqsVEMey7+ZcRvjwdkodpT89ivlKfh0kyLwhoUM8p8Ffpfmhd7/6pppe7oUCU40/zZfj
bkjzKl9axt06KXdCqwHGv5+plVZRthqQdKvhx84kdKc2w4z5CkvdIeRAcIi22aksJAWhq8DG4x5R
c4/Y7OZ9anfHgMiXwGT4n0VnfdNPw4fW+TiOG9aCIAlsOQpttRe4z9jOKNEo+b1RQFPHoP6hNQqr
gTDDMBkup2VRku0Pxt48HH/CXLS6OzQWTC2sIYE39e1cb2bAedhR0jyhHe0u2E3P+EyZR80A+t5v
/xwIxbJX0yqdpvW1XrgODQgxxTU7k4pwVOwKqSAy15H7Q+78mCYQBd6wK2vXBjIPXz+I6CGDC344
4Bo/ocfir8sUgXZ8ng1w9uqZRsPcbdStzppCSf674lovr3+204lzldVxGAs/5mjZe5K8+MtyGbPC
JSnt//uEyuxALjAWwR8o2j6Ct3BvNPdVpNLn0g3K8zy+1kZu3fykKY94Ql6FocBq7cvN4Jv81+Xv
OJ6rKXnQ+Jy140Du246XWglr443XtwQmtAdVtKMBYEHC54Jw6npq/zIVFvf4JIPadRMzZcDz2s2E
uiUPuETrN1ChCPEL/WCfng0RP8XSqinXMVDF2n3XSDPlEOUs5I2dAvn90848zn83wP8pd3r2dz9J
5tB5MggNe/iSFEOjTDbsKMoYEvDEaKBU9dkMxsQgKprmrYvesceVwKwuateRjdMsvGmtPGoVO1um
sp2/OvDwCX9p5vtYy8n4hYkbUC/DuUb/28Lxt4EjszXxgVwbz6CVBtLmLP2f4rjWPHzcf1SKQU0M
OmaImb6EHW4lqx/ZA4aSUCDncA+yFx3VIWI7eGSr9QM5W/p+8c1ewc/EvIYCNsy4r9BKvndlv94J
LXnuoMT8r/KyPfOYbelqQDffrkP9qCUv5ljr9H+Ph55/DQ5SzpCSdPSYfjmtTiUcr2zjIxkvBiTv
3fDbkP9JtTbTF4SLfuOq2UMhDxgEOgEnC3NcEg4+bDePhd87P4QQc/WL6kRmB0pHgUEpMHe+/ACF
GvlcIuMTsAzP1uLQWhYdVITE87P1RaepQFDzi9ssN+XJRE3HLJ+AE2ru3hbZmw0Lq43yH9KuetmL
gzjMhTHHnXGoclhh9ne0PE/ytRUkbs8yI/gKwL4r6rmsz0IPcSXOh0vg0YQ8flT+u0FA5//xs7kO
wIWEIKnFTV7zmy2VzBrXxFzD/Wf4mYEj4ycPl735BYazhc4XvP+4v2+hwzYpx1hlk1ijMHD3tjJf
CbBx7myT0eOu+xnrJUfjFQzr+nlGzBcIKGIOn4nt8pke8gp7nuQ6/c6ita7IoSRfjCLgiiVaLFnt
tVm6j3Lc6xoIb9bamTBYbeAkv7m6xPZ/QXCQwFlm3yPFfxz2HTvXwO+BlPbxaTTmclZpfW5tlcQE
SbcVXWGAftNUs8EgvrZka/EqN++OwNTkge0SbsOy9fH202sJCyC9wZbxCOyNBHi1BnbLLJrBaNCl
EHLrfPL+WOZB8EYvSlpWSk4c0nTdWgQgGKQdAxbzGVxfD3PxVfLCQ0BqN7V3ZESejRyF5XAd0BAp
hH9amftuZ7OsL/eYWFbR1BqkRKd9Jma94QG3TXxn4gQmg0m55M4kK51jR3nL4GFUGR5zLVfq7FNg
84WfNh+I2X/BzVCP9T8lhRaOIlLd2/KYLBZV5+xy2Q1drFqpS+xX7WKmcNsL4m9sGfUmCTqwVsZx
gGod9NO6r6lmhA0Ff0mAurVGYr97kXLaR1VRl4Iu5siWF3nGYGXC40ZsTTGlKL9mWYG6PXdYW2z8
bNnOubVOKS0DNIuX87Vn9maRcrTDQHaJe3rXS26H6gNvHHqLlfNh/e2cb/06aLQu+UudgU1huR8Q
/9RJ5xlvyUE/qBDMKnQg7/LOuRpTw/sI7WRigfhgZDllbREmctwY00uWb0CZo2ZGp6Cs/qKAz3q7
K0BB8+UUuZo+hCx4girw9BMsdxpEobPmoQIfuGMGc7oI7Kj/7U0oKEXyPcB1qlrAiTQA6X/tMLN8
D5lj6oDCNm0Tu1lKge8O4PYiWbGPB7/3D+LaBnNfgDc1SOIZIjKENJgByFQQEVx+VqVlc169QcR0
WmTiV8ULoWCOOET3RpXjQSwmr1E73NwmBsY0LojLIet1nSmWsjIaAtCB1s8d0d3GWjyF8FtDKx+7
jCorMFRs/Ah1RoQxAOe61BClFAKhUQg0Z/00hLi9cyAZnRXy9TBlmIbv9Bf4P9vMfr/Ua6beS/Ck
eHNGycHkG5jmFMdg4Ik7fgUQjFJ0rWpuB3BR7LOxaIuvOZtJ+38zeSfT9a71SW8JCcR+qZkoeEAH
vCNDVoiAYJ2OvNLTWAk9K7eVE0OciNDh4Fhf5ZnIRcyB2Kqam3w47X3OAAJIUyNXVpyEgM62vEws
0+pBLOnR9wpUQpmORCr5Wp/5IJKk7Fu/YFyw5crq1RmE7DtSNQBq/+EgvaSxTUoKZvhiWYdIPTG/
lZeIKeC6dkQAaZWyCB5XoxPYztirltPYvu/kuy2Uqyt0qaU++xUmE8lb7p+ZFs/L4ai8KZ5AwaJG
HcWXGuBDNxJu8tvT6AiJQ+MixjnsaJErPcc7uaLFPjO2K853thwRVo3EPW/lUKUyWNxqsK36c6eS
RUIrr2nRzGuheMtMbiDTs6g+ySxUjuVqMCZCZCxtBvOIcu8hwf7Cfqap7I+Arfphrf0/lhIjxsR0
amhKiVFBv3IdPg521iGbwFkJ96vmU7ZNLLhcrM5euYOFpVmlBRWjgNj45Qg7K3Ovk+GCA8feLYh1
GvUYFs2s9/X90fYlIdygNrWKUnIEjbeNglN7fBrztJp0EGXZeWlr41aqFo9Ee4WqpBnjpVgepy4F
F+8/Wh3GyfG9q7V1hOgJkQ3Z8nt5F9/OAtwUnpgrYTSSTFnBeoUnQCMU80ZOulGJrBQ7mmNV39I9
3hjT2TBoSqfxkne9N5WM7tgpYb/EeKbK/Kcfn43xJhW88lSmpWf2WtSEf3sGyyqzh3nvU6PxNwRD
ONd14Lbvu1TXmbM5HGYTfRWp2ALOn39mJilgfezsE7ypGwa06zVxdm8fiN8M1BAJodzhlKYGXgEj
vWAQZfIu2bbytWwBGncYlsJ8Q2M8sWqdacevaBIu9i8upoyWz0XCxwqhIQyUK0FMxGeUpPT6Xo/3
sEBu0fpjf3jNc3Fm3wou+J4itCUpyWnqhHUBTyNLmVrOj1saX7i2gi5F92bpkm0kpd2jbeWiZiaX
vLtL1QAxthGs4zZ19nr4anIofkjIPIlsukr8ukiUPJUbUpSzSBgniK4rFBjZQLJENMrFisnfluGE
eOcnQ/o3l0x7BJIUQUYXFaNKUVFiPH6iTa9Ga/QJUa2+uZjOAPvYC+4/vW0Ztqz8b1m74iWX8AhH
solEtiv3gG0zcMaAyl2Lxtr1bWFs64uhHh2loGESn7RRwoNjM04Ro1hZi2KtphgtOk3FNJpDnfe0
k90uNNGAUItU6imQ5o65gzDEIEefbDkJv7Lx/4mxjIULAwDJNFkB9qnfOB6DctXQ3mX31Z/eDP1B
OVpTnIXbR4jibqCUap0UMQ0pXEbZvzwno4EpDbeQbRAHlZg59xsaTrvHQXvoyIUsClCgTDuPaILO
jQO5wz99oj43P6sxKCak9+pWPnFUn6Ggt61n/IStn1n46ciLZc9Q4zwHgsO+WUXcDDdtGekQkLGQ
FKtpidQLJpGKsvRzJoqP5LZPJ6SYMgIyAX84tnA7jC5j00Rr/Mxonz9drDTVpf5mIowkSVpK9hLh
ATzlAzCwZWsOrxLUg4Ktlgvu/k5Op8hDIhf0P1LSGPUhBOOZhr3bw6WsGEPNmobvpFGyBCZO0AhJ
kLdg/kB6Xa2mXUR/U1Q8b1zkJc69ViPYPo43WFWYUaVzbPoim+mBmcIkAI6cBsij4bc5MJ40DQLt
Q0LCEsJyuuST2M9elD7zrr6PlrD142yPltMCn0WKeeKLq/FkbacIFSTqoCpunPCN2ZKd6OvGz20h
lpNbN585yj5zJisE6Ps+CzvCkMNqGz8o+Wwo2BjuwYJp14nXqgDxrPTtEZ7+LCy5h6Od3v9EOxBr
11Qr7K8Zlaw0fvGVWXwsHPl1YaOH1nkoAOlLhXVxMo+xAP4kfMfEfPYlmW1WAhVYvuh5SXKqiV8t
acpaRh5r6lKVy9PvM/Vh9DMjiufTs2iHtXNxKE4/PFstgencwZn4uA6K1sflPxDI3PGeGSZ68GQW
49s7/aSG7W7qfAJHI9z1o3eIx8AQFwaOE2kHsuLS/0M2Ud7btIEiUrZqmpBCYkDRYpta5Kb/6HFg
7CRnYJQBkm9QIOHTTME5afamj6aqEu2KIy7Q1Und91rNKenlzxNNlDOvl+/a+CFHgkaRtOrxp4K6
83I+3uM1Q+wTkz1GPFUPfZxghSqvkqneZ649J9IVywbnJyNAX4jYUHAc4NnyTKr21maD4NXFDpiD
kwDwHHLkB19SEdg12MerGVPiFvEW9xwrb6dGV1W+hzGyOKKHRCYeSXMNz/KQhtGh2OVUY1mEeC8K
oN4ej051p2kB9ka0+IFZWMNx37vnTRuduTMPTWvUMwYRVMhWHP0mSMXA5Dl7lEHZkdYqydkDaWFY
1ksDOQCfFHSBbgYZMJO/SUYgHwtGHs946jatx9lf/FbyHtLXisiDBKcv1nhRrm6xPmrn+mApku8/
Deh+59itJxfuwREB0ZnLpvLzMDjFBhbbZIiQmx9jkiZuIOb0UdYRnFWVEMEKPqLQHEviU/DtuVvK
NBxhnp/fuXowRL1Hh6R9nlq1khKHWslg4VPLYxVknOe55jDk7vBLGuWqG5ajZELZW0nuYDob1Qxf
satFeZ1yW0IyyqTrwqW1+3ihxd0e5MXMx0E0VYVryenwAiGUJQHRDMjt6q+6wau+yLy2yYPitY7E
0tSvKVu9bzF3j3QYRnhAWCKYmK98IF5KWyEVViPdpM5tOafgKN0H5AlbopNWjXTghqI1tcnfr5rd
USrRTpERFTaLA3mub416Ze3xa2i/VNLXkQEPeocV5WcUGsojIB2FF/JqEZ8Q/tl1d82zvzAkP6OR
SUZkyUgZdxLzXr1TTrJZwa01LeHHb7SIyZW/VsC7ZJYutwE2mwi0VNkhfhEkqly+9jn0DQbuxOko
uXazdmR0FRIbsC0NrpQyyG7gp3hDUUItJ/SW2oYsX+Zy2/5JxKam/hThBI6kYksbD2jXrHTQAMQE
KYENeVxfyQzFQvgkeYVAwUp61dQWjCCLU+RYW2a13+QHnTbnA8jwUDPKdHJ7lkkMCaT0QQi4qjCZ
N8+x4a0PCKNlkA7VZ9rL4uG2IahtUy80WB6asUimxs0YnaqtR1ntBp5C/TYWvJd4+v1ip+HWJeT7
PfBYWMNsfZ2IoVv/Je3xOin03vNtu0sE/Qp/OUyyc/UssK1tJfvzlowhJjArxgumWM+pSntDuxzB
58m3NUpJJ5If93k/7vkwfPZkfrwATWOJn93XOUftIb4jCZsDcaUUmUxgKieFLvXNXHWFiBnj9aqg
F/A80PbPq35U7h7Tu2jYJJsjOLOj6VjVgPUWwjFQ5RCJy6HFlQeJDePdcOKVnEHAjgWd/ZosYWYH
8jG8odZu8BKiO/6ms7gSb2+L3xb5edjyD9rVkHpsmirXH5Kk3OuuEsGP+DryEEUC19yYBPZchXoc
AFXC2bnsuV/tICJ6j+HpXE31xTv6PkH39EB8wVFHaG4kxC4VaPlZ169TlH482TDyDLQqS0buRQK1
iIl+LZwH8l/Bsu89qO+3YslF2Bis8HbVTlCyGaSe0ZliJ/9GXre9td1MYQineuG41c1vs7zP7zqd
ALEF6Ph//bSBvShf7GGAOcZJDf0svT3Rm5N4IQobwlKwk3eQ/ldKbGufF6blZbvAzMWCIBSp7cdT
S/6PAShrMNYv66Hi7jABUAVpelK9DplDAMBfd1uLRcjOhJ+7XK/w0vopQlA0jzbR4WAuQHPrLbDr
MVmqsr7g+fRQCbJJYZ2+eZMIiNtQqyM1i4oDGjsUMvg5LNJFBodKn8KObxLdqyhr6Ep5JERXJNX5
bz+KpB4mBbo++6MnlV61qtjL4b0cshhvgxOTVxESbuekMLwKQWt4i+v0nX7NiBOqX2q6Pv3DW8cY
felrMw207WlXfhNXbxOWV9ww7rYXpMINkq9yHWEb+FSx0j6Qq1EJ21KiayRGs2M6hMG2bS59t9IJ
57CEM+EfR8B57aeFsRRcKPxtw0IbOo62f7ipmQf/ZEiMQqR20kKpzIFKFTglgqMugQxP5EwuXMb6
oFnBqi3qkffM0pSCGSy4+kdSKGxyr4RGwUCFc+ID7mO13/22RWTQK6dNtU0zG7p2kdtqgbYkFEIV
mzvEaNqlwUxMAUDOx6pMeC15izQK3kG1Ml0YPVqSCQhWRGAUVBjgGJElNN+gYrjvRQSi/8XX3+HZ
8JUDvA7XH35unAbYlrqtF85uONXcVLsad7WVczVO191Ohd5yE2DO2+iqDQ3BT0TUMEIrL433ia77
ayM7Lt3HFMco/cpGyI41JsIAcxAynCa0itwNG4JsxfTekaK4YIOGTooibveaHRvrEjCh6XgH5O+/
OQ0smsHwP4YMnpJsb3pVOF+hMVxo5PUm4/vta1GQ8/LvUL0ocR4ymOfKDjmJhWRe54PLfb3kXjQ9
BzKJ2Mw2uNng7aZIZomYIFeRagbd4VsB7MX9YDF7aP1Fg63su1QK6FtOq5GLSajRzZ9reNqPZkY0
h9k8KiEBL6HxfMJGk2QhumJIzsePwdaK1/wAge+dg2WYZjWROGlZIr1TzIBnezjuSYQaGkxI/5Ir
35WPF3m11I2dIm6pB4bU1Vlwjet7Zx4JPrAznHz+ZpjHAiTvRrEWgRfxm59iODaf+8m9sOJd6JqH
WevUemFXn50hlGuEfOdtbJ0urvMx22pA5A+2o+yiSIdWRbIIKs+yi1UfcCL8E8WM4IRNJpkWjl2r
TmXpVGMnmexWcmiY4hJqbS9wOQRiSe25wMUm8VjLlAChfFTeXBXIlCtoxInYu2MxYqDMyALu6B6e
eVtZoLargg62wI8GHaHZqKiAuRELoiIfFRhAE9gRlaffN/fhbdijXF+CdyOEUmpukQW22TQpc9tP
xgE9mYGFcgI4CQ15OZoU8XuYaMsnCBAdAXdoEYGUfku2RowGUbN3vHGzyyPJ+FRqrWAp8JLELuVI
Z/c1f/8uKgsBo25txG1WSvQbDHtXZfSQnN3EZ5jnq/ojcnAtnoZjZL5GxGcp92Yl+MOEdYc4b324
FehgKa1WftPybxWJ2QxBbNN1IWcIEopkni99lY0i6SGvUU6BcSzSnafGP7TmjrdWzKjKbJ8JDIqw
pNo9VzSyyEuiQ/HtOYqTtwpt+OZ4LXNV1pOKynBQDzj5n6I6hwCGRYasIcp06TaP41WshaLdBXRx
9hXKK+D1pJvUkxtd6p+gszHGIg4sq5tTJDMk2XdGE9EDas4xlV/diqGYXMW0Nnjca0JVikeu8FOV
1Eis7zF78qIHgT+s59JQAsrz/8zpm5MrPIpcWqjrAmZCD1/gNKfJqR9KRPUCGtMDWepqBXuZmZgL
Xc6khyixbuFAlRro0dDKOl3+l9LJBCOC4qOfdN+CUqme86rCEwrK+/5/0/HaqajCBqIREIKQ6G+C
K2XsY1QNq5/tmflcZD1WZlc7GU9MhWuUqOJ9EQqiKOH9etTr/iCSJafmvHZppLIyebDOxyUR6KvW
S56XIWreGXV3S2ga+VmX2w9l/4OZkoMk5i128jkvWMuN6zJ/5c4kG6Nc3e0DMbFzAl+GxgCAwfZF
jDlz57at1StvTVX9CsRDbCvI4U+0tO5X5vycX9toHgJweOhtqL+6MOP7ui3d/p0zq/0gPP1wd0IK
dOxN0eNnD3mYPQ2AdDkGbm6eQ4ZeHcPnkX41PLLh0CIei+F80pXDQO4KdoUVa3YUN+1y5NVHeny8
xWEyrhGN+70T/SE4gXSnvQxg2IPFci8OjaT1t9PcRoMA8Tk52rxPmshJtNpdkRdM1UINKbhS+51S
IrMSuwc8QYdfIPrB3+Lo/7+DmmQ/Io/u0aQF3fOGXuTEZGmgQkdkZlVn6AdyviSGPbHSSok/PptK
Xk3jUmgQ/d0l3Av3NoxIgNoSowMwWQekGNojdpV3AtnfopDXVHngAJkaXTckuQlWglVD8ZlEeItU
okS6AOIWz7ZbPLiuMpZtZWtStSgpRIMr5m1SNf6XERXuXssCNDTy1vu6b7kXcxIq4CwXpS74RWkY
sTVlDeGAMI80t8fzO8GQ+esP/HQlYcOJrC4/52sQKiWfYwG9F6DQ6z1BYQ+5Yh1HoOH7caQ120Ph
QDgePYBqu9Yrb8Q57WFr4FnjZDN3zUqD86xtCCkoeDXPpjjR/gmla3Q9NIB4in2QTohR2/JAm6Jh
JLLH0uKp/yMq+GrSsp/NaoytuC+7MWJsUZCnnZZLi6j7j6RRDhcDuKBNefSLjNTYsXgy1AZ+eLKG
rUf5/JjF62l5d3N10HU8mdiANnINEQqzjDW9QN4jMyrwKIssAyKfFiIKOpE/esxP6+hnLlCx8VnJ
fdJM1XCW81EI64yFWDWJxHGUePRekXuQGzGn/hrIDqEWHUc/A4HBEYZcwJ1FwtOq8osj4c95pWC8
Jb+yw9iVsDWUPKRt+CYTfgOfyvTP1RrSKRwcACkBxKVsrj0Fty7u4Vop2yI+RTaiO3hpp17U/z5r
+bejLlGcPlaWPzH1ETdCTQE0Hvr7m8Jl2OGHzb2PealgxZnlBb5IwKcMKprkzc8Pn3sRXfZQk30/
KtcvnhbcAFcPnK+YsMm9dYXUM6GENrOPTc1U6nolj0sOvMyga9ngtIDdJn/KOo3xL93plRiKk3Io
+um0ZEfKM7fitLfTi8rbANuKYbOs/hqRZNm+y3A6QSvthSNYq9qHmB5Kx0lKyMIx8fDV4WTmpb1f
1euzq1RwhDeMFrCHTBqByeRz0FDXq4zDfJ5QODagga7wegbDCTVwiPRAHPruroaqs+wS4VAm5WCj
MWnhXSMPWVQ4hau+D2hd8U8V7r/iKleNfNWbvkpT5wtFOqBs6lYEsaGWyZlcKEbc696Bcjw4bMCr
Rze5diggR6ukJpQE1DFT4vsToSnheydmHcId/1Z2RdYm2C8rQ8PwvaO9GZ4Lq+FzDGW3xxmp8Eje
+XrqCBsPanKGQmq0MnO6ft+Tutn1oKOq1EGd8AoWmAyenfjHHnHR7UjQ6FI6OJLJrZyjAE7ROYJs
1F1PHeLPFyJZUuDZ77uo7sbQzR8RkAcvDnS/JYFIb/wrrow8N2Yljjc2wDUScBvDNlceSiPJgxUC
sJ1A+UCUJVOh4owptoGdS0KF6O+F0H83bXvuzmM0hVY7pjsI+HFeagGcLDFgzY/TLcesJD6coUEA
alZgeOtdOmqfjqfeDnUF2fwqEzIZ3uDGpXIwbfPKMzre+Sif66rVf2/B8Es96fsXtmbBzmyVLU57
tll6kKiobIWbd8ADnoq+OnDpDRhW0ZtMZvuQE3bDwkBQaZ9Nwc3uMeO97kSh6Flax1bQStaJefLX
V56+yKrMp7EqmuqZVY3JWSnGc1U4STSXBT2TbdLES+2MTJCM55GtmKDBn84agAbUdLRZ5arznIbU
+PQRuDHTrw8stI6iIp0C2cN/h0+c3VH23DB6wOXxysn+pSI3s+H0eoqlkDjamgBM8dqK1VcqzhLH
r85fIAa5pwArsb1r6WIZj+U0WCl8yAQJ7h09Del0gpRz0YCqVDyvVceGkvWqw+q0RtYMoUt4nGxU
wMngRAqt1oLsxPrQWb+jPskcrioH/Lg/45d0i21OuDA1v6bP2J3vjrSmM11P7VpfQAhJhZnyeMCv
4EV51B3NF3g6L4Ja6uzPgmbFJK3rFFAqeagr+cwqRgt6B7S8zAK7V5TZwtltr2hkQ1+MVuG9Qssg
DeUUEolpI70w834XqdVvxahewI8Pfa7XskaS/iDgKJMaCao+zgIe9KtQsVsawawWnvP77iQPnf5q
lFxzH715snCeDldxNW7yp/qkDuEP8ri+q+IOOwtoN1wx2xR1EL07zTeUP0By2yPSritqHOkVEKZv
Fy7ocnGxSDv34cW8lbzB/dWI1Op12nZou/IlsJ2cnf1Pi93F2ErzJ2Ki0L9EP4nWguGqDx3K2tAu
zRQNt8VCvhRMF+OHubJImKJU16GKMyHDquKPj5zXySjKh/X6HRWD9+M1h+hmz6KMLUnzTSv6zxzC
LG9rrung+o4rzSdXOnhsePZX+V9GGdQ3fiRprmWl0EtDwGohH+tkNPrdH4ewEtamHhntYzCPmZWY
cYHmcVmKRpxePPaTUhU7i17CcVqDu5za+ENldoM8qVMjz5ghr8KnGJrnPIzT/5HsEZFpYWTQ3iWB
cc1WHfTHSb3Yr6CNYfi80mlQ5283q4VhefLrUCcr9+XxDnLwV8tlk7E5MBQjlPhvwygfUAxcyTGb
+DXTXX2mvIZuYXJVMwA37RGgnwmi1zYzI/Cx/Of+BrGUr4jzrt+XKcb8pL1S2/TC+kItVuZcRSOQ
qnnSZQwJmy8/OYsc+sAzTuKKDjuXQGKpd2toiJZ5mdCQ/2yf3l9EbxmCrJZw9W8A9oiG/CO4n88O
SblkEuhdtQN+uCC01ugR1FGQRlzsUHUiT2Hhf7zIIWLQtSq9LYIiNNstRei8nfMNOTOu8IreWfip
JWp3T04UfiDjxesOKOKyt/FgY9AsK4TdnDLynbNaNF5XWAtJcDnBXuuU0RMbggW7Zk17Uowfe5kQ
pA2vHZaYRa8sBcH5uZRHdPpOEA/KLOtyXZ+kW8ScwwalgDFWhAfDm1ksh63ksVAYHXoq6cRX150b
yU4LEUED2VJ6bR9V8WlbmSuCZYwjSb54GIe0/uGLb2PaW5JHj+4svAZGTwFWq4nb3NxFDGnUp8GA
wZfKym/8LAe12LeLHX0vZPwHHPdXlCSF+GqicGwOuuCJj5XmGFbdQFIzRvQKbrl2Lg/ZxSc1rIsh
0a2Duq4S1IdHoIX3OdEYFJktvo25DjloD91P5dk9uDQcRW8W1MgJOc6/kasgbJUrSgB7FooVzq+i
ABS4mCLPQl/BzqM9oj6cFdW1XKdJM3N9J/k1odcY2vYL3ukqa0FvbGSI/uP03+1bSz6YfPCJjkzM
e9tHyIV5OnOi+8Lkvws8e+tMUMBHjybrUaAjpBkoiw9lip2HsawZ5LCfVdHT8f7vuJpMtJx20VXP
ssMKIswMgTtVyxLiF9fWOKXiDc6M5YjW+AZQg31wI78P4CHpCXj0Ggd1kwEvJE9OOiFtTMm+1us7
VuFsaU861y0uhoDId2mKggkD69xidyHO0oLYfUnCDoaUzTVEXGjUtgNBaRmldQUtzsRkVgEI6IPn
IIlTDfWzTeDDt4cru06IG7dFl35JzinFMAd7/mIGCIZ9U0Leh6Yw5SUb/kqJhqSFAtQgDWeh820c
Qe8PRXg5Id/0cUIlQCBmxdQQFLrlKUROd6G08F1iaKHEQV1BnyLVe8fcGRNSmCvFr4jtcQAmY3XG
aJVv0je4pCDtOezC8OgcfYaFIcDQ5D5BNLazZ7yPrV9gdH9gF8I7iLPxTqG5xzKfcHqDZhZGgdIr
eRxSjbYy6v6wCfwRyI8f+KoKCNAys+RAGSfOA2S5Xd4o5lpKrl+2ODkhzCbHC46iMgAtACT7nbcg
bnm8JpCm2P04OnWK/HKZVl6ahNAaUlCOkO/v54dQMolkzwce3E8O2qpqB5fg/lH78qtIiNrn6cfV
2CBkXfEpmnspzeWTHLLH2SwsuaQa7gdeDU3wqAKEBZ68VGO23MULQM7gzvwwHll65A24MO2Y9iva
S0bnYs9PCw1vMfqTjZKtDEt9tRVTTEyt914BlTuJViaxoa5dqBkCSKyKOt4j5J9IQIwyb2g5QMa9
QiYI/Qiq384r8IqQBeVUiFssUTMlCMbcXmxUqjfcHNJqyOYw9RsJxoFFepfzxhop9q5yK4jxqK9t
ujQu7zUJcGoqxI+h55kxrU6McUBocyMWDsUfEIGoLBVtjjMl+MCVm4zC+vicTQRyc1zRXf1KTf/R
3QBIqC0r2FZlq5bf3ZX2wXxSLDVaH55te95n6gW8A4JXT0HfnsZZ2C5V55RXc0mwc06QMgmW3YDG
SITOmHJEZ59bqFfq5cb/XaTVQSEti+CPBZuArbZR53AM8Acff/Q238AGLsRPbLBkw6nBPEKiPSDX
Bn8ujPtCP1UyHPic9/wgE+P8kEqHKlUZh7jLLmvIM4JHLQUKI9ooCcBNdOO43TIWys93CepdJClV
OEMYp6HV+dlzmW8Ey+a9UuqqtvxIMuOl8/Xd+rl9sMS+V1fjoeCIh7+sifVuuw8ZPeHvAXATMJ0E
U23hr+qN/Z51Frhm0w0apodi9Jq5XuQJewDpZWXqq/AF7NPbjfL6hhRGBQjr5C8r3Gh7mePqY1nu
XNZrdJjfVstsBEF7A6b+kgVJaYWHHGTmEJeaX7hwkkXJ28ijooMh27bqy2m5lA+OcH2Brg6PI4PH
UeeZU2wZGhIWDHPceSIpjf9G6w7yCdh/p2OEDDB+ogW8NtrXeWt9feoa6Bo+IO9nVrkXfePZXh9L
sCBYSf5af/6vo8kmNRgkVpLOQ0qL1Zd+acGsygnrQFeGedYKeT757nbmiBc6qbwsStYBtpL1eRrc
D/ePvmtLTTPeK+IapUIfHKhbgOtDNlyo8GgX3cP8/PiUj4gXMpdbkRgGzLzro5MDdmFGRE1CJvfr
nDQ0BSEORfsNeJ8jREiLpzkiX6nE2ji605RD6Z8ioSFUUQJpXqIMYBQnMeUt1hOSZN72UNUMtmQx
6ec+VliKsVi/B6m1cOBrBsgeGHxCLIkIa8Nku0tUQxCXY613E+2PVw5tZKa84hdkh2fSf9pQyi+K
ZbykV6fVzex7PfPSZ8Lmic4YRl6CnQELMxQl
`pragma protect end_protected

