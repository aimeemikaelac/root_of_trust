

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
cWdhJVBBx0U/HbQaUw4wfu1vmK1MfdYuuHme7o0Vt6a/IxaOXYdyrxs9okLeT3tslWSJXYdmqmDn
ZLYh7+ocVA==


`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
M4oYAM1DzlhtuwkxWmKCfjwxDC+bTPY55j0PA+EhnyetF1CdODudJt2IxI3ImMOzuAM0VIwOLNbK
jMC92fP2YQ8j7QBQkmu05UUZTePbshTT5K1/BGkoSAoCpL6BEDjmO6vq145BRr0zns48HUH0YrRp
jdZgXZDOdMH05IanEco=


`pragma protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KvMEG+F+RYYtbsJpF+u7hUFVxBvlypwoUJQPhPfb6rViAa7vM6rGxIp+X55NIMHhKYC2l5RZLLOt
ZzaEv8Ynprl6UWZvsw51UhjI0wWvw1KwD7M9us8QjbuP0OEOSDIZ1rpoFKmeZDT750mRpowsFDp7
Jx9QPU0KJcSSWIOwVeA=


`pragma protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
1osqEMEn/R/bha9mTK2Hcz/1PqMTn9v/LLSO6kyTXNqhmsdGSPiGuuKJdOCO86//GdF5YfrB/hib
kUisqYAbHTAJR/bZjxqU6VOZHtY+lJuY7SLT8uiWkvtLeFpLuIbceeOdbx8sRlGXrq1nUpsddAZN
Vu/J2nTML3160LM06f4ipwiZBD0B0byxubUhAB47WF+KHiu/SAjoUl0eo8r2t1hklTcuFe2dxtSt
o3Gz6jX3iua7z3GfGsGMHzdf/8n2Ioa51ZXfo0HxWt9JcgtEu8PlqtGdXjuWU3xDBN/qLl+U8nnO
orfQXhw0wSxEtU4Q+6T04sGBXBOejycpboG7Pw==


`pragma protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
piclQgL+98nVOBn/u/pIauk6pHC6ljQw1eOi7JwIzoJMey4lvWMMbscdNSVaxFunh/W9tCM2hUfD
+a+C4yTISyM9RDrzHS6W7azooXRqiSnGjBQgQKveZCWbUY8J2admgWVTrSyXkPt1zIfzaxXeY6+M
hCWXWlL85N0TGRyFukgWiDHEiadBoqWEXP9PYrNSkSJaggxTYOzOz4kthy3JuP97HT6ugXo5d632
2mIo8Mq0PJuTbRFzkSNug01Boszfm1qJYwKJfYeO5A6GrV5xQxOeuhuQdj5uabez7G+IXL97PZ+l
pO1iTjOaPULSSXvYz/bNnwORe6XtbGIhHqaQLg==


`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
sTd6lvG+mmEgYUbvXuqZYudrLgxIw1ZGZbJG1rq7nV2ZigScIjiAxvliKfLEDvn94ki2OqkrYB6O
Atyx4FfSd1zuItLDYff2MXkAMzZR8PNjNI1wTKhac6nYbLZn3kfGdXRD8FxD1tJPrve6LnsXNO8r
mUgJhBum2kE3Xcj9wqbwesI5r6+s8pkaMh6tD8Vmlg1WrUXhZZHZccUtVhGPfJPsJ+7irG6f+nu5
dnzxQNMNRFKyGUOf1yz3QHlqAa7e+FyBTL4gKezMhqVkzOpJ10XYj7sXlo8lBf3auXfb9Ne3hFua
LQx6ctTtYkjfmYnUae1fN2/I1dsICzB2JXjvBg==


`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 405360)
`pragma protect data_block
8SAZ3OwDekqJaQ/g6ySv+SsG+a73UVdv2VC/N+1WUU3BQQri1JDLmj4VmH1+p3GEwBYdAMrs0O39
K1BjIX3rL27p3kdWlc8fRcrAi75Phvv5pQEU1Wow5FhmutOsOeTCwM/5bq7dGlSSNQ3etoi+ztdg
aeGmBu0UHzV5JaErZunI6ZGV35rANpIf6CAZnn7YFTrbF1LZ9moA2wGrtntiBZoQI0xSPg+SDgZH
H6KKxhCg0kbJ5ExyOm2i68CddUC91XdnW0stUurLJSD0yZTSLdy3cBhf1vDE+aiKQVj4pS1bCBw1
q4nLTjdQulASkPcab+TyGDvNpzkwzmybqUIkLr6NmnGj+4BRKAuv8Z7/ZSGS9D66ujzy+d6daPZO
1GVfyR16Cl2K7pRKOgawoTsKxldstZRbU2NSV16AEAxlttAvjWU9qrMr6qy8YWQrXj1B4VqAG30p
TUyxGzFPTl3rrXuN4UxJY6LI1BFhhDcclfOu7jbtC3J2Q+jQ8FzYN6HbqGDXiv0e3qFpTaumaqre
vvVRDiD54cZAJzn6CB6KtaXlH1lXqQwpKTFRIen27qOfZ0kATI3wljka4nh/3drzllM3BHPyzcmn
t0BtEAnsNlZSnfPmjuYjDQl3IUTcSeIAlp9U71ExArxEbEEDz37RfRazLaRRRx/NU1TBtJEaER/f
lvjs08T06RvQ6V3lslRWjTXUKvZFvFK1t0tQ83bOTqOxeZQT+/aO3s/BYsa61AWH9CTwbiar5NOV
OKzpDxjyxKTCVy4QTCGX3QmjVG1B7N24aJVJodqEC7osHAtkviSFV7pY4vI6FPmkPy/rUd/aR7ef
09hPA+hUryTEDo2srhJA5CBrGg8lQgZWHozWs8eVR3GLug2iL+1PmvP1cauVc/mdye60OrT/htFq
P10Sb32upf6qx53UJvdXkkKF8FqhieMEc8MQfqhIgXoM5lE3jMVgspbTRThvsaNOPxHJ06YjX3fr
vWJSTQCW6YlcZAA8kLqwjuMCPTBX/DuvDAABn0ocWj/ZUKaFQ24i/VeOhjfu1iPL7te6vAU2RxUi
DByVk48vW2fiNXSK2Ce9WV5cB5LBMbWtf6dfJ0M3dCxNGbabeBkNbJDNnMnBW++Bt2/wnHs6Ckra
HzJq3XdRB4t3cddVc1OXHnVluGPWNiUaoh9UJ4cvoeXU7vm8xAtG/NIb+36MHI10RIGUTLYxJwuG
PYbza6GJs3rySCG0VXOWubGVOLVk49hhes/Tkzl7CxWgYzco6HJTnLhVMBF7mIJc8D53+czPS2sr
oOMKzvciaDhlNzCJ+nmFhAbHuo1WqpgX3Mc8w08W9SYRXzq2WCjnekwPN+xnFwyS4JyWngc0pDDx
qHx/Lnu1MLG6Erd4oi4QXSF0y7ZOzYfj4QOctUKfELduXeg/ZjtgaQGe5hSMyK0fhjkCSqT5lbXw
6PyRqwelKg5u91FbAF3q/ekKs9YKVEgVihw4FQTqQ8fyO6sSxxmePa7Hgt51RlYOHQAactB5fcKq
At2YseE+w53I5pwoZWiGMkxDwk9J5/+XoyvYSpe9VSXZu8zBVCHSIvKMvTmXhllPauBwmZQXrI34
F+zWNoWns6eQv52Jf973vtWE3meguWfEBDA6eHwoyM9DiJx7eeYTHsYgZDWahKvRT+F96XP7PPdZ
VSBKXGCEeNNsPps4YDDHxOpX3+uouTCgX2NXtaT/lWYYc5GcFfYIM62QNPfl6HqD32fbGrDoJf2E
8brXUA0XvbGlhr5ZN4/WV6MHqDQnvMrEGdZ2P+tJ+YRWXq+0d8ND+ga/0r42Torw/XJ9DmE3mp/0
0ALZ8BnUB+rRzEZqKDVSymvkjH2etQ7w/MN1ZPAY2g2YIlAtsTrqIjMPmPa/kYkE8Iz2JfhcYr8w
6elINRimmqxq2OuoMKYZoKjm5OCjQpjb98E3jN7xtfTj9CFvcRZPHpkHGKusoZaSTbFDn3ImEm6L
GIlCc1e8YHxMG6kbvueZreGKnHoffmYcOpiAlu9TvOVjjQkVMkZV8V0ZWImYui69IFGap7KMJnSk
okXoUEy6Yf4vXHuL9unQ7x6V59dU+DeD7RjGwbvxfaMXOkOp6isAUqKh4qIkOg4cCy2LTeT5Cc0Y
PhBeiblLCIxxAzGX8X0qHkfdFkEXVBCOrwBqN4jKRkTd8zgz1A8+kvPsgwuiQMkkDNrMuCX+lBXg
ZyDnTHINHNmzo8nxByH8Z+KHpzhB+naK5hIFRvMCgZ3+qe0g43p7EXBpc+unmqzgpO9nVkEMdNmK
F8fpa/UXa2NmGzTLt96zlbiNj4fXqRwVVpx4QIP2pb3FaakGCiMtzTQvMXHBUxdArnakxIehVIp6
fgpsWC67Z8fRjfXTvjPUjvvRrThlfvggMalMdv/p9hGVCApUKrxbPd4R8/wqJs7ctpq6GmZvxiZn
CIF1MFS/2wZRu4dtoMt0heLDngkfn3Mi5MIe7LMXlBy5EZsWKyztD5dTxjMSBNSegRy5JqfCwjfv
ixVwgeIB5FlVQZB/VheWRPepOAnV7+iDMIuIXuKTwwXmal8zog2m+kIbNM9SK2E0rgM5w/Sexxmf
86bxsMitcvtfkDmv7wMQsfn+8MZM7RfgacsAv8xWWlQWDNCU9S9pkIv1JLIOxX75phV9tn4yRPPh
asdD0jdzL+YKZlMnB2BfHLYthkkyNwaNmQ15emLUelg5LMc1wyhyGGkLaifOcbPAURv81Adq9UVi
bBcmgiGCiZP/rk3Yr2aoLRDvnBnV7sJJgDHZXYoYx41edBah+yg8ps0vpYStYJM6YTfSYrQkD1wy
XGkHB+LHILPKg0I1in/pJLUP//gzvONcaPssyFbj/zvqnTsJN4znAYSuCaO5HNc4GyS8qslpP2c9
TRVLJaYzQjMGzheKAAVKxpkMd+fqHH2zdnsvDSdeLPX7hJSwRo+lkxUSPbBJ4izqbUVHMRdHV0dO
B311cTWLkvOyGwIjGnfqtN4gFQACY5tkfwWOIl5hyVo4iqg/tC1ihF5goT+1HlJdvOFU0MFZ03ZN
nInDy1Cnr4uh8hLgj9jwYJakpiNlLKkwfjC14JT58+Toua7Megps9wM8gBv8grasHhlOKXJHImyS
fTDbpCeKjbcGAOBNxfpu6LSdeIkbBOuMzAnaQRP0XuY3Pvzrhqi726RsLv7n+yOPIuekxHSbhu5z
ilq2DqKxkAavfT3VWhaDF2xmKiJ0wfxURAXfv/onWdHO4VxKJdFogML2RfqKX4F/cMyFC8mvtUYM
6ahn8QzKBPIYwvdP3Pjwrpy/4Fo48LTb05HcXgwMUF5dy/vcmBrXuCFP8ojOP0CgUedH7d2AdcbV
n9uwo3s81gxABe+wt6pXVq60h/mhVqSjrtT/39s2dO6xTk21lZ8EjurCsBy+4QQui/isdo4NrYYO
CP2tRW5f6jBSjUISobmV7IAiBOVy+0QfgvOIfgLLc3p3yBO9ooLPDLn9ffJJIkbilL80jqpUbQ9L
ene64O1peBFlv/NdzzoRQW2zTob4OupAE6AwMmAI1XG1p0TUOtFiWwcuzuQZkF9o0oR6Ciaq0o//
W09kc4wVXgYbpn4RR51j5VjIRZ0kHWb/3rqk6YTSTCKUrJZA8I9NsQ0JuiN2TValnJZlUR+lbR6X
TxU9FcqcDojjbEJrNuYlHO5XEgOxcT5bxZJTebJ962ueeTEiyYnRIv4chDEn1vkL+Br6BNQ305n/
XBBRY2l0M9iY+KMoFrL7zqVPATDehKNIrUXMf9/ZKZjLls5Sxn7IvZd/AIQ2gE/q8e8v3shOQCRG
/fU9al/GtY1DgICpU34kwcoa/4SF70zNChus9AFYW707ORsAZa1FB6fffr4hMV8gIAHgJgtk42yD
159MlqOB1K5xslNvKC53b/DwEIG0jETKDbYNi4/4+skh6gXkLdPW8hjcRx57UK1fHjCC3BEl4Vus
g+Q577VPwRkiYaZ+Gua7QmvByZo46zKaffSPtaRfdVXs6ADRMEnnsbHHuHp+20PAMhfYRSf9svRa
d37x6VZU6qFODkjpIMvKVf4tE5ZAOQleic2PxtshkvETymxeVau8aDCuQBLd6qpr1wsfyBxbIOdm
j38P1OsQEEIHQbJx8AYVi+jxCNJ6LSZPx0tqfCkPCLIzowUiPmbihqbBa+TZFHzyuiNAykW06ndJ
2vkGcgJGRQApHBhYrbysfxQt+1jhZCrM5NhDDcnARj/PxtoEsogakoGXUjFt84INuDpITCH+JCy6
Z0hJ1vueNWZR2tGlr744qT/SsHlgB+w79ZVGhZWqEx5HgVdUlvZkDccbNlExOlqme8OprrSCdTYP
x7ioKGygp4PACuEccDTBdTm4j1wFiLnfIQ19CT//g8hWyaD5NDmV7FAe6vNXmhtmj7o/JWE2yG+4
FSxZSHhboI2E8jVvj+C85tIVDNhbLVgz0X0MU3Hj4Igs9RxhwIGkzYrz9GiBSeXZzy5qQNq/rX0k
5SDzphS0aqPKDwdKYyMEmHxxPdblBah2g0zH4toOC2un4uhYaCcMUvyvd/0sSAIxAH03ca/sehTF
sPLVHHIPxlyt+M/V0rFG4mI7zVVt3iP+qay7462gt2AG8CbbR5NrNhBoI8K6MHnuA50ZKopm91O6
gsUyzi7FgYBwRKGHNnAYrhavsW+Bdo7LDim3V7dUb1Jt75lKXrIBM+mou9wW+ybMeuWtkI3BQE1s
iXH5G4FZu7GOpD1uyF80q2/YMivXFH68vNnsAH0gtbc/V/vZEym5BD/cCrZRgacDB/9oEDZTJjF8
3UjovV0umyferX6i0VxraQRxHGtUtuYVIvgf6ArG7apwzysMIFtUq52OI9YRrt/HDCVCyVrXVGxD
GD1RHsFgbgkv8qpII+RSJBCnZpvXCqG1Sbs4Jc/G97+Mngf6H/ltzNjAsdDNXB2Os8SWiFpA1eP7
pyMDzT+Qlvie8Mre2MtoLQvutKKksMuDqIpHjAzVfcTmENPtxOWVd7MDMvyJGaom4pw05jDXkk8e
GZUYnyt8v5sxNDyvufeK5EngkrSBJ1t4+XBQ7SsMdNH7xakKjYCComOOYPaN1kcRnpZokItrj8C3
IoZmm524jsrmHzqikTOpswQCVCV0BzF2NmS38nZ3SOwiqPH2fZoTyTay9MCQW9Ub2mqTyel2p7LS
YbHTX5znYQBJAyxTYnATXInfTCF3VGFD/gIOGfqEOzflkUvV9vJ2q2ORYCJ2gBq24/q4+m5ULvHt
cXbb9i4YMFd9wv8F0XNmojygIXWEN+9HwJb5u++K9AP1dU/DQfE5QSERilEkw1i+dy2inE3C/qNw
MoH5hdzGjgOUrdA4EMuLP+x2vXxeenOdXV3C7QhXmOWGM7MRJhkgExC/KawFO1mv54LYnFoCBIGX
H9mR58aRRFu3I6wZ32U/A7ZMO6uuTc/2Yp0TIlMub7ogHVOA9SXL8ML1NwwcP1RVy+WXDDIowBuh
gTdnBAWQRqzZwTDA8DFLO39XTH9aqE57Oxib/xDQdJH2A/JFnAeRrh2cQpwIv5bF/1u/h+p5Hx2H
vrRK2qKXaB/5Pu0e/mWkEy0BL+D62RbMro+lJxAn/sBfh6gakdeyR7cfTyxMcOhlimPlHFT5jT9w
BHDqg5oDun81D0FUh4xP7yrId/GwiJCSfSKX95hLoZ08zSHCZkXmHB52hl2M3g+p7GKZBT7r3Tf7
epTCWuxP1FCFYe7CDG9eJlxc/FcVLw6m5jGY3hmtSEzo/QML4nBiNnWNCXnA5+Mfv24KBti6lphD
WbNu+tJkUCZ1iQ31F4qiUU5b4wj/FD0mHyhgQ+4hFlihCWzVPM5KUzx4XB+TBikfWG8J1/rW7/Xa
0VdCkVyxRIRTB5YuDYOHRAY0kMS/mLhk6tlSXKGBtHtnBIQkZq1yJJ9Th/ZWDerTaoTQmHM/KRk5
Xce1A2s39H17q7/lGJAyUyQt2Eh2aFd4XzAnjWnv3/ZVH0+NixUSvUHLpmq9NrIQBc664zZDNpJh
8gFY2nYwv3jvOPjcwEA7jz2l5tPsOTbFkT7FEdG2clo1vg2vmJsjCNY+vBGtS7o9j4ZP5FJ3JyXZ
VjyKpZVQmPgHnV1gs6yZMHIsA3auW4JRetcmNUjPDeeBBrKkKXm6wQ5nJNlKCwVK0F+3f7nIZp3M
KlU5JwzjA2aWIqrpdMQdyiL/GSvecTw2OpXApQte2EBgNQT8Q0YfTpgBOzxB6NZ+WsUTRWZRmVqX
gDVCwPzhjlOaDnY0XRpTIBRKqh7HMFyUUesm8GQX1Cx9w8Gty7m5D4j/pHaKCkNDw3XS9edIw+cM
cRz9mkbyUrg4VklsAGMRENHYQr+CpmPjRo5YMZQkKONISHWmr31rQGo9wK3UWNX31DY75wgphMPd
GE6VeKHviwcGVWTlCmU/Iw0T03AcdUUM3biXneFr8GDBk2YgOCOu5+cKrTzo8PzfkQmEG75Mbl4e
4L2Fk3Km2CmuO33aFxksAAr+w9si81SRJrLilRrfIs/Mshh7fD2jUvIP6ZqxhfGM1IXyuepQxWIs
Z8OFrEAPiFD28/V3DulG1EDOAEnZz/akHLv8KZ9RKkJLS5K2xRmnC8YCPb/i6JoUZfyeOvCUT6TN
qfA+RPfIHui94n78O50VFJ+pi+62w9kGB8CPGIS2hbqTNvZCBJ6qZNygH62O8yQhVQSsbS7bag0U
zAK+0zqKkvoljZNIRWgSaBsjvs3gfo+bM2n/2zV2tJSXynelfbZ5d4MG0kN4kig8k/s31a3XsX+v
1b1KXmq6+Gh4UTuvdWDl7MKX0zODJ5x+hb/e9yOBuzg8Pdabg3P/7nQSNnpHWPV52KCefqvDPJkn
qdAFhSSmmJGcddrxTaPJ5OZUVggulzfauVTYZHD7vGmqtb31qVxNv+dVf1owfQEUfFI7NrCXFvbq
XywMpLZNJNDUzexykteM1jfg2LXP4wuF2GeaUdUPUhDtAd3TDVDNliZ2M4LmRZyQHoxV16EYnJZ4
xmDGcHzurx7tS5SVeuFILomPaxR0lzJxkNbr0jK6BSgyOg6l0wa4txtwF0JEK0r8Jz7YR8Vk7SML
h56bz04GJxXfglQ++h/C5lWfRaNe2NmsJiSHhHymKWesTniAphtvpqaQPMwwxMlbQHrKla+vcyzF
BTPMeqZ4CT9gBgbh9e1Yjy+mPjqyXHUmKRxyvciSLxgxNElq+jxJ2WoL09s1bkQpEuwC4xzF0Cla
WNDy+7l6HyDv7mXoMYZzgPNuvMO406TnYTQfvEof/VQxfQWTG57DhlRbMdtLv+ag/hzIV3sBt4pK
7xhFaJL4BzwR6dpA7NdbZU1OAfLQe4msOzI4Gt6DIHjDTJTyE58gNqVhfRk0938HJKzj3YrwgDXl
FB6FSdYGK+MPZl8gN/nUVPtrImDFdBfLveADmTjaF1OyTeMSnql5mgimTtJ3y+LBEhsmIh6QsqaJ
FjK7CXWNOhbj1YjQHDywvX/d2IHQRQHgfckopJ+l8gxGxluvdbwNIFHcXhoH0TGxho7im824XXbu
NvCOPgv+F7ER5J16RE0Bmo3wuw937+LvZspm+MqDghoR0icFQAuNfNZ9pm9cNNwtj8KfKwP/0z1R
EixG+5ge+QKq8nvxnNz7WHpLlNIgPRgZyLq/1tP4hHIGjawYvhfH2dMrcavs8HuJELSUkIRMht9U
fYWGGYBRDTMmtIfuQalr4OSsdTwYysktS4AT9dlKJYdqJhV+Hdw5wHSsgfn1f6frba0d5cAz+ghl
tmrsDtGM1coV3e0zp9mYfj9UHcKmAnObU/v+21O/yDP/r36Q4GTpXGtxaRYwPSV5SWPhp3fKAh5Z
yxsoKd2t3JecxO/iQI04sbnxAPgEGAPQLvzoAAboIzvoLx4hZDtXVPv1xeCi/EjHWGqO5B4u2cy3
8W/fPaSc/c9VmN09VysOa7SHagqhtXTGfhYIkTujUsJXA//I2/iIl8l8D/RD/v3v+jILN88+6UAU
9uLFZ2KAQc4Ll6eYH6rVnSJz/hfh4g0NX3rPMwrjmap0PqQqQx8MaUqEGCrUzdJ/6l+X80RW+Wg5
WNaeosht7on4xnr1W0X3Me6h/J5rZl35z8XEMJSNO0yrhdhyNODlUBXbtWbQZvLtDEUlJ2ZQ9DMf
IYZyA4hl8N0IO7/P9ohnwVbSLi9dGcNkU87tmFuytIw/Q5nXZScXVEmjDTE7BVqjT2jbZ3JXCOLz
2qSsDvCdF3Maawdzsmt5l3GtqCKBPDND3aLIrJ9exPLPqmhdK4Wd+VYOX5l2kHFZcPWQ8W3Rq1z2
EUX7ta1s4nTlI5Dwlaj8A3EzVRZkBLlKneZuGfqm0hFWcp5xtmhXACYkOaKqsfW3+NX4lfxgxCn4
coE/T3E2LADri0SseZG2K6CrXaqtynUDyNZobnev2hXRHYXS0rmtlJ4cOpQzGNEr2gEIEXezdMYc
1E67LWVOfz8aPiFiS9R+AzmUnjUBPFIjNKP/0zCVuc6t3pNmLtHWIXRfGBEjl8EIrbnGtsZk94V6
21tidBeuWc1JzZcGmVDbBghXJYpN/+JENx8+Mk5RKBS5lWWv3NMnUlQqPh7kNzOVuAUJ9/FjGrKg
4ICbj5gqIQtFfUV3AasUMwF7scqx56s6/RZm4MSLRa2fMeRmi/BwxSQm1O52P738qAZx29eni+wU
4sBzxtybAhlsfq/PFO3RRByde8eMWpNA6HipJ48ow/HDIIP6JH1wQf0IFWr/fLtqFScvs1eFSrqw
y6LJN0KBCIUPfPQivAu+O4Q4lHOBOzISZW3yMzL1uvGsZes38bAqtG/AuVmRnubzP8h31itHvLU1
e8m7u8q2tM/3inwsGUlq95JadHTa7xvHCTc8C1daTQQkVzE2/dzCbQQbl83bjkPQMGB3fIlZT1nH
ZOktc7Nva4EBU2IdcHyTOTW5iMGRJlrd7zeOAh2YACp3EkYAmIwLQ6zYmvBSDuOmmUMg9TYf2/g7
wdLXY3PHbdZbL+uzvqYPzb80pWYgymP2Fw0PlvQJixXATglmOsyE9IIesYR1gxcTy/Av19UQutJq
vAHoqHG8W4fYTRppIjJ0FQhwTwBxQro7NcXIvaryptBvJlzNo7nvOaIrJJiSiEvfqXS+wlN/tX3Q
8fg8qOQ6pWIhyDo0OSN6En2sx8YhGKe41uP4cGNFwl1RuGERumqGoeOwYmSCIPx/HPlhyKECGjF4
iSKtKfraviUmISRrji5CzAR0vbj//TMP0ZruP3gvQafdY+qwDS3TqKdNOsYDMh23j5g4NGsc8w0a
yclCmUvgp7VCwN/rJ5QSlwwGpDw7jSgkFInzHy8czyxw39Njk/hYSXnXDeKje7b11ig+TO9qtnN7
7QHRMlOc2svWYBp6+UuVSJxWC7ew2N/F18A+vqFCQXBi5Tq+u2DkUvDZ7Wcm3zf/nslAx3vcxppz
MdKqxa7Crs//Eroowd+S2oNirnUUtgaU7kyRXItRub06wrtM5IBbhMZbL/y55KzkWuey6VHLAW2C
Ju2Nmw36+4wreDFtKUWkRQ+CdhED4ehmVnBqXhK1/eS4WyV38DJONN+jWjgFAr3sbttVAJBttoQ2
OvfGvZUK8Z66zw+3QvObNOmxhf4dIQu3/vFX4ti+BjElQq/vH3utFLE8XVtmjgYr23H5oVvb7eJt
D4GtQubw2nE8/2hXlbHEejLhbY3GgLFSI22e6WDUEvxbso73bdu8X33nz8j0/71U6YCky3A6IYPC
+KBqGyPmvfgCLZXwQ06j9pWycNlDWl9minkjJUWp6ypEUuL2oX3iPsgDQWPU95Pf0zKTk62L6XOO
j/GoVu/WMV91nAhsK+o169AysOhC4YXlsxQ8gKLycTJa+zNRNjR05883bIUWxt92A8S7B7MzQL31
o8JqN22wPxnvFeAnG832hnNfT4jTMSx4CN205g5DYqxZYLRVy9K5umSKxegnrziXQqtLnQSUCq/t
hocUz9niqtmumvZL1kZs7kyoW6z67xAxcFoCiHS+qH+Wa+lOL+Q44M7R0DC0wIx70ssmtILIpeI4
ig+9fOVlFEFnsSaqa4asSq3jkyl6j7CSj0m/avooCOgtEQ1o41bow6vcGn4HbqfKDoBTiCwTcpUg
HnV/c1myXlTz67LapRJ7hCnAAeF6k/gXQIhNbCKIFu642SF5ZAgXnpOUmNztAPdYJUbR+2H1sjsn
7o16jMiQcddcCPe3WqNI6cww+l//YU2XJuvOl00FLCKHj8DelY6hxEC2NgP/pG3XnsaLwUmOikZh
+ic3C6+H17ppa5BiZWePHTpM1Ga6N1g7FGscWBG88u4f2lcsidRFYyZ0LFRNpnibH0BQuq/jU2fq
j+061lqSM0fZm4pTGfG6mxcpx+TmvoEY4EstV5G0huj30Gz+dsFZR48DPVWLSuzV1UmM/4NPXvMV
ZrkSLkbWQuwjwwfDw1hF3lI+0rYSzk92O9Clz+FyLFWMK14+/ysg882KVhqeWpKJtxiW2mqP8rme
Mr7pnmZnjLlGyh3+8FsVItP95vYtcGz0NuPvSZq6/DhyTI5jXLgYQvMOUXKh0FCnyyqsPXFMwsca
fD+SINQxGfm/2Frt5yydcoEi5+uyl94Udulk4Ce56ARUHaFvjmMId/HmHFFuAFkJNGaD/VfNtuj+
Ez+rvHVjCalx5PbOTDqUS5sVUNHG6HRdB7RWFjfaMZO1uK/dLNfZErLQqip9MfP3sQaUpjR6pM7K
lQRNTL9q99mTWkw/acvSDiM8pi2fcANHeIuJsAydWdD4vnXquz+gyec6s5hPeoXhebBahJ/6hiaV
AN73W4w6jY98IxvcEmVH9iwdO0+LeAnGOyvzQg7eDwWj5p23hcwOokVRrC2fpXBhdh6WzBgWqoH/
cxTPYghHzdJn1oQ+RYnNDYDMycEMWCfnDoTM1I7OWElN5h/An2YFbtDYR2ukY42vYYaDxm329ZAv
mejlfhZNHfu2ARReaSXRMKmOJw921YtPV0ABGaPQyemIfy8KiZ6vAlDFhRxR8/p7nAp94ntxA5Sd
gH4NbH6buO28osyH2h0cOorWipyJenCwr5nLbNNMFJsCypSmALHkYdWDMRz1ASIb2HFYdoms5Pgh
40JK95UPr1eBrbnw/VMeHZszt9efn9rY15vINLJBmsn9jUOpoiM2WjSIOz0f4WEyzcTYz+TWJthd
Pf9NGLOndnHXl3a2Js38orGKn7CsORdvdlDYi0pdXc2Aguf2Z5FseFtpxWSaRFOPOO2zdP3Ylmqd
QvFRs1Qfjf6CW/sQBxAYwW5Fq3w8Al4Oxlu/d0xmcDprrhPNxOFAhwYO/TExXPeFztuxBX+GfDiJ
HRfMua4HjjezDdg+xWcbMVl4GOJhfJBOgtHPV8/AoRKiufNl/gjbq331KCYsSr032qvnL+pB+WFl
UKK7ggN57oQQkFVrtPEiIXT8Z6LbVs/wTGzub2s7adCT5cQ1TvDATZSRrS8SMA6R6c5JsloeSKaD
8r/w6L9porwdLzLYfpmlJjzMad7ETKn2Ikc5yBcCa4nDNDXqysEBJIOXF7/Whmjk+MfXXH8yw1h5
Um0peYaZTMHM6p0LT4CVqsIzD/nAAOTQx2F6P/TvTsoEMtHjfcsMP/5bh/4LODqpsFX3H/9R0Tu9
7OXd4wlJ/u03jEORA9wSJh9C/0/EO1oIr42pgpzsoZJrK76FhVgem7bOBEiOA/u+hmOFRAMhWVPa
LNH86xln6wvKdmOOJk/A17QPtr5Bphdo0urT2TTQyCdFgBjr3ngDqP3k6rQ+MiXMxIFqyzgpLmTu
lxul1DP7MubM04hEH6k8LdFIlc0HIVIxQbQHxAGVR7uybgsBPCFQOh/Bg3JH7eDZX6PBUTI6g+LZ
ayOo9JSANoZtiBruxuNUH2oTWV0mkKQAiEVrYrxd7P5pF1N4y4WQ5jj+NZnsNGJNf/0MUx1N4rZw
iKCBzz3/WS4JMYZfXAAPIBb9Eh7n0ETwVZ2FMUtiKkhuTAEnKtlblS5XCBseZMJ0jLItObTsVDQb
qGnqIHirPCG/VaGP3yWBDiX/qrMe8hlGpqpVMm6WWiQFS/WODd+iSWP0S0hXRN5LNNzgkeIROOYi
LA8zC6MRxY7Sr8shgHy51XGoFxw27iq7pAMKz6bjDDadWNIkfDyp226qJt0vV2wh6r+QrkA6lrOJ
fcoJ51LPHqOLFsuVWaDklgxq/4ivKfNBGdgqYmvn+TkvXDcMJrhy5Fk8RRTEKq4zSngrutGNKyRZ
6UvML2AFBriRhV8Aad1GWysGdg1iziP5ZPVdctklgVXurKJAAdxJLDo3xOcEcJ0XJgRbrkBj7Qjb
KyjuLeOciFeuATZMXxtsVkwb3/Cjr0hs3b0VFryT2/oTQ0oZqev0uAu1xgzR0rW6xX4S0J7fD9WI
w9gzX8cHXViMf9j7Dz/ZZUGTkoeIZPsGz7l2DgT20c8R17vKzNvc8HUpycAKn6t/KyjRPbbnZI+F
bolYVBmRl2E2ZEZtdbDN4WMzz4N5sbGJFUDIDfvYxmALGRnK2JCmgYti9v10IOc7DT83p7CS/WtR
JYp7D7Cmoaqu2ZUoheyfGMwUbjBnKVonchamZqbY4fiW9BbEWPTlCLBntqYmctDaVRcnsPULzM5H
uNqmnJ2IXbyhkgnM1VAN/cIB96JH/9TSroWDRVmSfojDeqwei74XbxYJYwXDkObLjJ81NUVIppQ6
QUAcUjXgbE3duF9kWrhi7qH2WGKk59bOZrhuVNhkLMFTQnKO31XaVw+8fZe4rM7Yr4xj/eQsfX0L
zoJ3jtFnJMtaHbbIsXHblitUItYdWI/6xEMxqrN2m2q83yi62eRBH9/rcK8YAjsNfaLhr114zaNV
0LyuTkBVVo38P+Rp6iGy+mC8JyEDPZGF75EPV3NN5MlvLSXa55cys7BQMMJwULi71cl16Jh1rL7J
JWjXX1qyUb1II3jCAl03Yo/PCByLyZr8cASwgYGt2rTKs3NW5ivEPPnrXurSrDpKXldvNdQh97+T
rLlQKyQHq2+6Yo0uRC8T4Zt8+b2RW3SCTrer6mmTYUFgt7PSEuuBNkZ6XdGgpB8+yuYceQgXpvqQ
BYj39wQkQxTk1MXOHMTwr0rloB+jmKquF/bij2jNwr9758x1sMdltPpUP6Gu9hOsp5YIyKJcp2gY
Ex8JfD3Um/4ehgVHXDoxSQpZRZRTaB7UdwsgXVI+eHxdEKxvHlCeIi68+pbNYLB9mF12f+Uz5FwD
TEVH+sEBF1WnuIiv0ZhmEa6DluLmS7bJpKQi8QHGnK0QnVsqnqTZLvz2r7hv276bHoQQa9NNCQss
3lGbFd5B79Yeta9V2iZ/Lc7sPAe9WbeiVcCHkEQ390VuZBSlSj6572nBt1dI1pbffvg88FkASmJh
l7mjggL6mJG4VNyif1sK8qHMywBZeinKUkEBNSdU94F/8al+BGCtGILxjnlUOxicNJe0HFDTolZZ
SnJfOSICE1XMTccEqlu4dhM73DIN+j7pElSSmobGyTYkZRxPrl97Nv38nAk54kqt5oJ2c1NDC+hc
VIY3elaZEWd47G3EpYC256nvk7KdXqeRlPWZrs1GGfdLluaioJtL1rL+L/YTASYkg235sHLTGRjD
j9aFho3r3JLPVONl+HvKB0RJ3teeyJAR3kLI/wi2nIdFLYQx+a+cMtUQeHLrCic/pC8Zq5O2pGok
i+2is1YYExJ2a8JWyExfH5qadkvybs5QpvMXg87K4Co+smXOIAOyBs5a5wu6zotSiz9SESHzD6Sh
+yM0o7/1sK78hBib4FvqjqbBzqA0eu7/YQkwsV4k3taxzYjSt4HLh0VRIKLqXRvpFCL3ktnHKevd
ZWZgtrqlSgXbuhaJ+xGdvLPxUdrHNT54joTfw5Bx1AhF61NkP4PU1X63mMkDfPe03iNF1OtVwg5j
74ss0AWSRtAJf7Wisnms6sZCuiW8fs62KI7cz4KJpn61n0QzkS0l4+vPDdzwi0ilE4wZpU34Lk9d
8+93wywa9qIEhABNcmhqTL01v0vOwNfR9wqpSWtambWX7X9ktPgKOqpIvZlvjFEgrUQcvCaDEX5o
bbT4ZbYJmwo/EhrUCR8mKjwa3+ZErTwxgcY94/N499CI8iZOLyQ2pIq9Wk5+bPaa6b1XO4EuFY0s
FfMla5SZxXBygmnPder5UIfSRu20g9dld54lx6gergcjlxjTtGWXkJQNXC0lnoA1jjnwFJCkEuPg
9Tggs4h5EpETimxstuS6/1iZkagp66iE22MawRFFEoD8mqFt117LY2/exrgWsi0GWtY7rRFt3tPI
XZgXmztViTmrfbDjJtZkjiz0uKmrzviZoCv8n/b5beCmOd8eD1jvKwD18wJZHxIPk+qH3UBefCQr
o190zKM3uiXg4ZoyLWXcKQX+o+5v5pjJQwdAnSyH1drWBnBQ7MO3DwcjA5jkvGKn5BVoaNUv0SLX
b+pJh3U9joqX+Ma7241amMD9IJnJXo1Wr0x8SN059zd1KL170bmWQNDCZsalRyI/RgxmDh6o+ob6
TUq9CdjVklqsqpETgKVFnnRmTJE6BxZ7BKmRaMiBkYXwqstwJyUmeqmONqWlaax9JgfJ5X2L8/aV
xDdWkp6DUmqLXb8d/C0vya7OmOWHxbuCRpRaHoDKjUzd0ReO0mPWsfu4dP6RbN5MBwUFRO12x7Uf
Mfp6yfRUni5qTs0RA+4tJSpJumD/xvHidQcpQ7MwzSlV+yEXYl9qZIcwxXChvo1fNHwodT8qF6iQ
tVqpwMolRrx47kdRld0aXeruQVZJTABeBnN6npP0n6NPOGIR1f+vWmwfZSKCnlsz0WMbuPrVyWXZ
wxRRFdRfoY1Qr1XIuB0QpVhfrs6UnjjRAp+MF2kln2ecP/2tjfK5thIFEmQnv8n22r0Fvs2iv38y
Y3WYnT1twy0w315jKWmGqNOud9q1H2KqoFfG9ZH1iNfp4oS5+IeH6wRvC5Lfyx6tifQVfIo8HLBC
PJj8PdrrmdR16P0xYuBlTgyCUl6nmdlAH+q3rkg+UM/aRDoB55fEVlNDMCAjMnpSa09eoVMrWbJ0
f54rqCJcvtnSokQM99uDCzkM//62gMtv/9wsXbkK775rO7alnmkIuSPKXdL0utH4kLN6YdiIoDyD
Z7AY6YRQGoY29OtoVKvfabOqvd9YPnXBbM1lDce9iEJ8g6vNqmQcMnY0cZ5/jjEHGP8Z1uTzaA1L
QKSmQgQg9jQ//HIIeVaarrBn5WiDcxVSA7Or1XhZvlPpCv8pWk4TS5BQvc6wNMhk6oA6utQxy65Z
5z/w8XhckdMlYY5b3lcLvrdc2OPhSfa7MKtYtBT/P/U9NyrB8Fe4skKa1IcFmfoUYtZMEtClUOOh
OmYo0mrMHM6UpBL7zwQbB0rM+xKYJCkY3tqN4AoQYaqjHVLS9tDLqx8i2DxA4vFUzSFeyXaeEN9/
JHA5X4uuK/kHEkNGsjg1y1OZNqoXXkzgy5hC/2HHGb9P/6sXHmltw0P+cF6N0FPX/dhBYWOXGsIH
I9lEkZs7uXKkj6eJ24Zyvdrgit9UvsUVvlkAKdJmfxGD6yr9cqUN2hYpEOQ9lk3O4c+Lq3TA8oxb
u1JSjwzytRyPSBBm59JV7E0tTsm6sDHuAgrZmvtdxoAVMkqBN3e7PPpBsh543YW0fWoMhrM3LA9r
O5Pl4fIC92DbB5kaKn+0h2biRi8jNN/HFlb46/BFIWbl+AFhJcNfXiJkMGXGUFZBgvRMEBvGFwKv
gaIlK3yjTw2WC3PChmsp81YUdr1bL1PiMEWBwGDBPO/IzSSsPcTLWRvEN8kKsWlgOeFNPvNtC7H3
DCXWcCJo2GgKWZnvgCP7ex+ZxC+EA1gd0vWJ92ZywsgnsCJ4Nv3qcWhRjsGYusD3fK9UxoTrps5U
FtVmqgwPiKHV3GZqfnI5pP3+xdP3+hORggC/uLjQtEsLzdbEtpRvS7SYHi2DqTp64uhaMabLkuyx
l+YHI0IloKmCjATdbcSnMcxV5Ke5jcc2SZ4nSmHgtk/XPzPQeSoQgU3HExKILm6x6/XXP48ZFD2O
uX7zefaF4Lve/uz2bI8LdoDmRmRlOwyi6s0xHSQP07/mc6TKEjO+FWtBiDqvsb9gewM5c5wczG91
bQS8w+yLzM6BZGjF3sMp9gcj3Y3whfJ/kuqUupblZX95B2xOlimXXDtI1SVhrPtsysAYL9a0e7vR
1Um2bgZbBZmzydUUIdcwB9BGRKWIS7U89abkQx4TSFKCJBXt5eRkwVR9gdr5F6CrZA3oSADx4kvT
xJLGPCNB5meSo8zp95e5OV+EMWsHcA5TzkfRpVbC+MWBBpqmWCWyYHGdEo4lrhKyxZYUQ6CqoD9e
7NHMvSULHziXJ0HvZxcwLgp7cSHifpxIwdsLnsdg1yZQ7iwWO6M6t3+yQDRNe+M8Bw2SCsjA7tzj
S7U4YP/EZVYAEUUs5PmQQ1xEkpliNW5JujdjgF02By9vOr7gtHcsoPpgOF6UyfnQcIdvXBL3cT7D
qLCk3ibZ4L6zRUbPr8sIViKk4w8B2GzBAXaPSV5LbC9hGQIIwz1XtQlaSfYhNy79tvIF9F0aZ3cZ
gmD9HO6N39NmXhjRqD5ERNnKkMGggg02jklMPSTOZqYChJVAkITUocI6OrN7o1r7ApeFyfclKU31
eooIkjgJCAFQqwUSViM0190DO8EdJIvAlqBpbyFd+h8xSOb+Rvx9BIt6vPM4sVomiJtZAqGO+2Y7
lAcLTIBNPuw+uZBeT0Va02IsbnMMULA6Dbt39GTwuBYgyzU81qoEUHISijFirb+IBisWqrgghBqS
9WPCTjC3rfjII11hvL9KaSXxEK3Y9GyLijnPXaRLobmYQpoyTuq1uswi+asxaKwv5su31iRCKd1T
K2KMLufeMoqPSNJSN6ZORGbIKIsYZBvd0CD5+UAihxk0g3ezOqO2c2C/CHS3LOla10Ly4srYq8yX
cGspN4viwXnEXonW1XW4PnaIqwDSrvUEdpsN1e8dsSgPiYtFN9DmlFWc72Cm+7u2ZsDFCi2LT7Ez
X7/CZrtIvXpBOYm3mJDvl4nyiYHfW6Yq65ScIdLjUl5WBg78MRoGBbzrprmpcE4Z+F4lQvjbL45X
dukZeYxKaPvJliIbWXxQeU6oNlIFlIr7XtQorYcYYGePzphVk+sIRGeGed9z+ih2BDMjxO9SSdfY
Q6sFWQzeSA767jO67H2Xrv7POvnCJ+YHuWeNtQZHVu8iBlL5/Ow80D3oU98XOsc+erz1S3LZsAZl
Mh9C+CBHEhV02LK5jDS4UmGQyT71raixD7BV+anHSrDgJl11Uo8Uh2C9VVwImbdcQs9CGPkAYbiU
14lyfPCuFaS19/7r5D/g3IhCiI26kg2sETeDbkG4IKgqE4BU4fxCmLerqpOWeSWzDefeFbPQpDS+
5H9eHRfm8rz4gbb8CUiia1q8bGz6tPjeQF3nzp4yPN/iyT0D32ganQNz6nCVjxwCILqhaC0tu56o
x2JwTt1H3haWkFLO/+OBxPSZkAVt8Tl5O6AZz7SE1FsIc1YPj7Cmf2GKRvC/8+1Y8ov90L/efgfk
5XpGOuou19m38+UXcLhCazSVDliJHDYDFZ9Qo7oDOKGebRwtLZyHuEjwhdVZ2FhvyyGek902bHLI
FNCGmtfyepNiJ04YEPPlHQSGC5nCY89pZPqfcScdRHe084NUbgjl028oLY1mBDKGOX5noSKSS+M8
DMANmkL7ERlt+sskiUSEfvIVLZoTfOAlOqOqE5NPrURsZ/9d0C1pU7blacEFuxYUPZIM19vuBdJv
gkTqWml1Q85/kh2Vh8MfCtkg9tI23stNCz+JL0EmAyjn6kSgPA+AzMUVM+hGTnypA70Nc/ADmxtO
hfLOU7MYvdfdnlo2jcgJ/j7L3INV1CSX+vmGj2f2QaXF7igogzuERh38/6MkYoSRLHumTWBdWski
3nmh7lB6heuVKY3A1ImSac3L2jJfVcDFHg6ae/EZKUDTHifTecN4sP5WPPSAYj8lgKaOb2h5L/32
UbaCQ7EwF5qoOKNSbcF4zb60aC38Ut9xqv5wWydyimnBPDMnFnY0yy1mIq1xaGqdC7DwzeO/V9/T
mYOL+sk4fC5BvkNiDbSv03IWw8vxFl+axG/m5BdfXPpAdqLRswvaDusLTPcbN2mgK6M/GEWK+k0z
yt0groUgD4l6SdaW1ihqcQ20g8nK1CknRUy/Twnmj6t+cL9sSTKLDz6vr4lIF2bQvjFKJuhvjuYU
fbOmNd0ltNovvQX+AJhoG+Ky7XW+95rDLDbujvEopmChEBlHr0m5W53rj9Ze8Meqpc8T6NRaNfYB
EdzKgzyLua3xJdrox8hmDQtT2Nlp/PHZFKuh6j37C+vEPuDvq2flCOR3nRj0ysviveLfIhgTUbWp
dBRYhljq9pjoCrOwebXkB6Vpx28nP/N7Ju4bq4CN8V8ND3QEzyoQmIagD4cOO4gWd/Hb/zyD4lIw
W7B4h381rzNJL8tahnar3CyaBovM4r0bj6jgYXIxUSYh8bwJYSlU2+5yRmLcRdNZx9e0fYIx/w2d
J3nQTqO28rChQ+i9tISqCJWrfgjImyzAp4wrzl4mKs93d/oWGf5cnBx+qDL3POSIt0BcexMeRXxi
2REH3/CEGdPBBICI8wXaIvsnoz9qJelNKhpcMsbdG4dfJNQt0zaU4dkqOB5ab6HQnmV3yH8st3Af
gSNgPsd9rhpPy6s9TJWGFI6cfYxtqzTXyao3IkBAedTG1GaBy9soMVM4ygiwxTdynOmwcWA+c2dW
Y0u2NvGKdJthOWXUi9pUkwdwdVQe8CqLTUZFAzfFialXV/9zLGnlkk1XuIzG5i3qg2z/RPr95nM3
zNzNpYb/e9SsQBKZEF/KDOeXuIgj5oh3ur+qWlpXP558AoJRK4LHsv9qUuEm1TNtjbEEVI4RhzCC
tJJDVnSMlSyR3IeE3H1OOPQZpz5CThQKJFS/o9shOJqVxHxjh/ietO8sAVDwqBbeak7kLsYAkoq9
utK2xwGZGWOiWXlosIJFejzYCBdCK7zLzduzg8dN+zd+9jtNOBl44uJKerOY5YQS3IAKJ2x3O072
sPK2HIAfR6QF/kdZGuY3LfwQuT9rRDzfX1O0XDwD+w19kneUm0SHdDY9hC7Ap1D5RFDZXFtKpnh8
3035AXsDE0hGbuCc9Avkb1beZjhM0QSqs0CiUBxrlE3hjSzdi2as7lrddp6ScFhkIvfMR+E4oRPq
BB+fWnyfL+HAjqQBpMKkMGad/o1RSOUbbjEDUYsVaclhDZOm4+DogeNA5xGs777dWNZhqqBsPDkk
MOzamKQUq+sfZO0ZZoVA9l/cYXpGxB9PyfUsPgZWXaYNXsYXdRuai8M6Z+J++1FO7hS8AEP2j1Ns
JMw7++f80KMtPF3N4Az90W19YYuzh3RmOQmpg55Zx7VelPGjj/WrVbjV0ThtAq43VeI2nw5TU1JI
dBXRg+sywTOMFehPOivd4IT/iw57Mk4ZKSqziebF+F08D52H11e0r5hc485fPkIAybClIWDdXz9x
MnyuB5oIY+BPW8tlWRssILiU72VNwkLO6SHx5Tc725gQ77xIzZu6AwlWuoR6WXPgL3upe+589qXw
KvVs6GR7rvfnhVYcvmHKtvFimSgvN4CztKFA1aRXDZuRjxeoZ5vOQDw8wQPVb+6k8GHDP0InwmKN
zYOpwvmNyD2skCCaB7QYjgIow+NZMT+UkmvOw6lFT69Jm45GkMus065GwPsBIFCd3C9SYdyipwH4
q/arBsnNzkwdNPX3hZMxKTgxvKtN5wLWGyu6dK5lZSsCg+nhGEdo6nEJHreLBgD0Fi7X8R3S955H
AIGlryZ2EP9D/tJ5ubxkejEiTtPEFAt3zIW9A/4S6yXnzaCnv8Ou6qqldiVXlwIw8rbD1SD7gQdM
Vip3GgjSibtKG3TCJmc70kNErZPyazHAYCgzTjoeHhZpWKe9hR2wrV6mSnPCdgI/K5bnC9KdlqB6
+olduTkm4nO7TKm77C21CTlINGh8NI5Cf9UcUeCa2IG1WTpStHBTFq/noWpIOEj/ntYE5/Zi3Y9A
KE6zchFe84RysJWNlEN8Y0BaBbFJwA+dcimuouwyzjIyqv1fNBHnGjlRm21AHKLO+t7yrPFkt0LQ
z8NYf4Onp5GEdNrba3ZD3WdW1Y+jRe9u9AyF/iOdo/dPezMdb0d5dCSpSP6BGU/NuRWLzScezBie
6wNxAZJ3JAQpWyRN/4gVrCK906Pqr3uYNem/zbcJSV3oOyDVKGMODeIpkSWP0Dy5wo4gHkiaLRoU
hc4VcqA+79kVNrGDU7EgTL865x5uNN8pWA7/ivSTpnOgeRyKZYKjL43rx6xA2PIFG0QDbkum8KxS
6BBJZjW62/HjUPmDENrSWndsHDt6orrDQJh4VDAl45hQ+qPNUG2NUNNlcQ6aHdqlAn24qB7tbSVN
CC5Q7bNx0//gZra4tivQ6dN8KXgTy1DjaWYWcNvX6HlG+/MxofuA59KafgvTHkWDe3Eh7WXwEw/0
DtyGlRm7HS4wB0U8T1RyBBDxQoc+4IzrKWiOca4Wt1dFPXSWHyxgYyfnGlIYtLI15difxIGrxouE
CA+IZ90ilvNMHPmQqn1B1J1iLvHZXvAUb9gGZhEgrgrcXkAjDZJ7i1Q2vjzDOPUxa6Cw4A6j2qx7
OPltd57OUBsyDkJOIBnEeNlvrrkwxCot9eTp5u72ZYxw/90eiFc5ip7dcNF+oYHCCsNSIOAGvqvC
LmWcQVX+NsdMFpmLCcY6eUNYkjH1cFcKFiI2ZUQLE2FzFH6w2wle/Foh4BG2Poi3YQ+yZbqsYzPT
47KKjvT8YK1JJAkuuZIS1eLmyTNaUq2HA0APuW5sUZZ72Fzslyrfrte01w8jGgEPP5yV+hXVEkCQ
KGLBdRfs7g9Opw2FKnxmB2/ViNANvQBce11x6LTLhz/kyDpvE7O330ValuSJZaZZzdRnWbpFB6LL
2tKkOA9TmcLNbAVi9ndAC0m+vhwEUsu5ZM9Q6qNstNyA9E0y+6BMdfvRY16/HpJua8WCpTVTtoX+
tKZigHzfjURQqPGDSVOBuhBVnPtH1nQSZDCJaOJqEwsPcgyP+FYKi2kZCwPe2GhG/oUtslPRamD9
dWsgNuZJxG3KCXSSAIvKr5UyADdaUEGxoCNoow31dAhT7AEwjiRTwxQBxodNYbTZfhxFZszmeegn
74o/XPg/TQjh74zPii8aUqLrvnEXF63WCJdAbdYOQ28QebatZnH/3PDNAazBipkut23awQoUd0Hd
YVdi9X+Rxqp8QB4bGygYkwAbangi7V1B1OmEABZFKHSU4l8U/jwhUdSUOo/y42tjBzLM7iOs8RO+
L29DUDbbYZcYq9jVIBoiL8uvc3D8t1k42BYCpYLGlm90WpcGyFTfOok6QANs6q1QkAlY0wvcODKo
9OKJhGiKqiq17CJ22Ze3kfAGlReOim6Nj4izQgSqkRQzFJhsUGyDMBa6lKG+GLnWXLYWXoMRtANL
d5rF1NILDo0EQMoNKFNcEULF4TDfDUriiXgWy7gyxhbLSK4B/bjEmXTGKCHE+DsyrBxro4xJ/Tut
SRp8Kp1l/g1g9M731udwp5oT0o+CyBt7X/WBmvcPf65W3GwDpD+yYs7hay3hP2KYkbZn0n1ItBqh
KKpFGcrtrLSv2e2CYdTQN/r1vju3zMe7Z55KK8ALC8mYprAwl4Gp7QAUwr1FHY0BhgIKd+pSDOI1
7NZusmsShJ6QX4JWrpEA5tMM6lg/e2pvlLy08EcAs7askuZjymg2oRO2yPXT4OOqfPJ0m6wMC45T
CAoMG2BZHmPX3T595iFsFyEQED7MacUZa+IqL4M2VbmVnn/Sygy1SR8UK4oaSgWcnDCNeONLt9BT
Mv3tNbAnplw8fXjFNVhzc6OB7zsUYMgemGvlMC0fKPhE6SSFUbMUvmO9Y0n1b50ueNlvfK31lwR/
haite0JRQFH6s7eegNI9+084quWHQPxy7Etl2vKu4OIEW02AP7SnCLpJ/fCfBDh+SGHr2ueiLy5n
aIYm1fbSPyPwfLXx9uKcsNHCm2l2m6y01e/Motip80vFKEQWp90YtDSPB0hOisVbRaJd31zjxIPD
H+8/PJZNDaafaUapCLeZC427y1GMYOlPLov/Xo4dtDuoBAgw42B4Zcoe2Z976osepahrE4FwqzJO
Yeh27O9z2Aex/HznKqY1BSxxz9yMdfRg6KrEk9LAxNwPqQmj0ow0wq8FaLoUpRUv4WO/2e4p69Q+
Nf/+Qt0vw7VrHbXzzijrGjzco1IID/zduxxgoQV/9haq+rp/HOkGl7rp6G/sbsgvCxzzsLPJCgxy
mxHZyqK97x1JvgZfjYbWFMuV/Dnz/6N2gOy3o2wvOcenK0CgOf1y9Oc+BVtnrMbdRfQQ27dFS2io
YJHqkJCjXEakUQ0SIApJ4n4bm66aXBBq3wuMf8OLSIJos/xOFReFPmTSpEeTlJ4ZxzkrSPKNnBeU
G0Rp7ZK63KyzixkEdH3Z9mPnv2dhNklDHBdMdj8l33d8IYUqKn8YY487C5y55n750RsSXUIpIytc
pmOJR67AJosfXqOzpkGyOgWTHNWl3X54fGjE0k3PNY0F8SWcR6ovxHss2vDdda2ZIa8Ci1uDDhK6
lmqo9wcJQyXPtp9BnjPtrANKuEA9zbc1xfQPuDblU0QuJpLkOw6g+rmbh6CcezMSjsoI9bUz4vxP
e6YFiwOvxYAdFhskIgvEjg37cIW3aoCifKg2dieobYGuiHK3RDe2n2gzehXrTH8BEJZsFwlvmh+L
nkf2uwSZPKhCrPvEPe+8IMCMxEwmQ0kjW4Xoq/Fm90aTsGvUxxurJ3gGADn1kd20ByunXxvrbbnm
hWoyxIpfbRYVu/9xdaXAPqOJ+eDTEkZyCH4c9iGh40yLDCKb1DNhe/gnrMFc2E5TbsHx4rpHKrHo
/BtpU0h/PJOlvvwW/+39RBtV2NJaQCGWFLQlQ1eqGGXXOhXk1AoGh4L5AHOxq7HC/XRTJQ9EvU+W
NZCYUT+DbY5iLn82bFY+6dtbfwaECoU/QmFOcrHsqw11tC8cvAB5Yq+fC5/DirKVQiIsw3PJGAE6
nXkZwzBWeM5kvURfWjQ57qSieD8GnoYBLX4E6vZ9aO6P/PjJFJoFUYJqNmrJPG4zYZV6O79RNLC9
K0WvaewdaTN/3kXdKbQTZVgbeQ4EE7+GULWSB3kzAokYan2Byj2cfiUajQJShf/nSBdpyBTQt5L2
APbkd9s+YfrJdx31VDjzRAua3qtBSTWDB9vmC1HaoCkJSRtwy8iAI8ipU7HofYHWrlHUY798eeSQ
QwoMqxj9i0qvfsDvQbdCHxhXsQ8wjR4Qybh/oznNmfcXXFkdtLg/TzPVzTG39Jh3JlkGgam4iStk
0qxRUrpXS2Lfn2sPa3MJlZ9Z4ULPPf66zcISvvIw8oCf0lxGNY05lGfScYRlJ/GsghQw6orzJ6vp
y5MAyEM8Ju/7dy1F7DnVIICeKJlj3wAEwVIgwd7NEWdqxoLX+Z3Fq4TzkQTkl8NS3Ir7fy1eOc+C
XwFmEokdY3CLaGb/+Uim4DSf2nFf2GzxuH3SRPQjrIAbrydG7+NDC/m0ixWlpG0yO6PrLvC1hJ0B
QLercLYTzaWvjoidWwOfltNlfUgcdHtrpypZxxHCNbhXAYW9bozYlgDcYRJ1hEmdeeDJTZFmD/qd
DPpblCwwbH+X1VrfBiXHE4lUD0zgg6mZKeLWmhs85MOaVZjkVBE2LdaO38n8Xj3UXHtq7AiDJxSJ
DzhG+SG6OC1M9tMgixAx8MjqUbLbgsbzuMsQ9sjVqpgKvQFHRXIeh42RjK7g3GSOmNYQKWY489/4
BU5h1/zdEIAZcopOHFyebRmjeU/BSkaSrac1idppbhwUwQtMupod1HrR0Yqrn8sacoG3Ci8GwjKE
hBFRFilJwJfx4aMli9gLM+i6RWs+BgQ1DKpAHeY1a4g+QfVgnf0r5hzjjdGt/1MqQjgyQPSFg71E
4SKdiwW0hlESzZ6+VPtaBYepCbpnjJPiaS02UAHM06noH9ZUFP94gWsWf3OVGvnWBtxZOlC5YIQY
CFq8dSawlSaJNwOeEziZMQ6EH3dRM+dJ28Uo1YUI5L4Eh57Dqf79Sl4UuMLvqObhyBEO6ATKny4o
ozx8ldWaSgIZohloISBpNMd0BtSsxSafan23MsfTc8FYkFALv4UybsnYc/yrj/9RA1lkI28lTuN+
8GRaTglpdQw8JwG9udR0NMSSMGXj+fU7j4wwQGqi33+aO8eQOAqEGvElYD2R2AlTVk+6Y8fGQb4f
O3ej8v/u6y80md5g3dKwc5dPVzJIdciebKI1cAJM+luRUZnX9RD+F1WMawbG9CW0ZrR47hw3a7o4
uEX2HFxT+H54zxVD/rwqRM5xh8q17ctL6Lpq66Pce3u66cmUD6J7fDHw9ZX3iEsKT8EvPAf9VyLv
p8dwpNYtO+5R3i8SJ0FvuLaDpWsioVwLbEeyi5qLC6nAaMFdc4xw+Pe73Uh1JUlyKS5AXebB+iSA
dTUd7JyfzYvD3B0CKNuMPGlz1LHqZxIp9sT3lbENMXWStRi6sRgW+LoqpBrQk2gMxLYHlyO39Nv6
R31RhcZNX2eayRElAmh5oOyejVpGIFHcvMCTXCL0J70A+uzAVQxRzr/5V3u1o0/wkpdl9DHqG9TG
qSFQPiUfdtZpn/0+AXfCn0C0s1qmaLqGBg3Y6I2MkcvrKbv6BP1BjwOmIsrmI8DyUYW4fc4z94mh
+SKN6DVUL32MCHhlClEcyH6RO9F5o6jL/4d40nQDuUuCnpgRYfWQ81F95wt7uybtm9MsbTbggkiF
sU1E6xuDhkQKrEs7JL8wTSCuMhdzGdaUilEUjnhYNL1RmrglygtnlWDRZ/dZFxsu5aZundsn7rsM
aQ+GS3pEgUFS9YyaCdx6v+8dgQ1C7ESoSvp3ypiQmshOI/+6wvk92r1qelOo8qLJv+JG1NpHzqlV
wjP+Zmeckp5PdlZLtlVSJ/IW7c5mW2eGhTVZzyrmYpOMiTm0MVqR3aYemZrF2LhvutRXZrurzO3B
YCQT4hStSj+tIcdooF0FSRseN++d2XCuXiPhokr9uW1qTLroKcS3L5NeHYeAXmWfEciPwjZBK5VR
nCYmvv3vF19NgSmShgM7KoWVq0TdbjEnolvmEvvwj7IBD2YimEDJ1LDZJMvTnCe1VmcpcVvZLUi3
pKSKhrv8YQIX1zkxt0NfGia0wXFVhPPtHztSBVFaEcEkAEiW6MLpNNGkYsetiUl0AxinNunSRwu3
pnYU7kNS/CgxvQZQeE5fcshBc5ugI3TfyPtPiFouHAW4ftLxgfritEwb7pj0wdyG9pYBtSCJRfsU
IDrOzKic1oBXLAs6K/+DExkxwS0vhWZbxDGuh0vuG3UD/2N1pKbnI3zmWSaFW8l9GBvH2feWpsCM
LQn6HY0j6rP34VsPgIgiPxPd5RF16Hfr2/gDGIQ5ujHquaroJQKAgPr/avb4g9wL9BnbKEV/3W+1
9UwS2qVBNLvwerHhzZsAi/aNLT9fiPUFYaiIgltEKV+FsqVe3B0t8sEn0mcMJQiIR9B9qFIEyDjS
pMP1UTpHAeWifEwWYrkT5i0w7jmNka3ot93o9ROTPVB/dfWdxC+VNZ2552I49+BqAiOE33Pqy4Eq
qheNBfYxtDlEKK9g67GrJfImw7cnCSRG49IGlc0CoQV4Gc1eTGRHHnY93LotpHJHJPysny0Aqlgd
Z8eWL6RhZWov01wzPT2c4SZmDwF6W0iqHT/7Owwqgo84uyLoBhodPaBURiJa3p28wN/KDBGQxyH/
G3vdoNZDyx8KpU+b4FfcMrVtvASf/WEwAG4Ojlz944PUQpwYxzKd+oAVIuDPJ5T0RdYndfYcWSKF
DAmyr0lh7vz1gMtkPa6nHdmGHrCqucsvdwSmDUIXe4ZTexFlIQrKZC+xfCBPkuSe/LdtjPoRCxK0
uNz/lZ3LNXGDN2rorA63AYr+JhbZKSaK6uei9QzH1hWQwCQp51j0KnF/tYNapjXxVMDWsU4F1mgR
rm7IBPI6o2p7ouVvw6gFQdNMbeXx1Aagtjnw/XNa72u/PwMrSIrdJgl3O1tiLpWJQbw5fd7vPNFk
FDz/lzS4dcqYBccaRh9NYoBF6zdHuaMoMl2k1ufKQDrLM8K8lB7UY3aJvJbQMFc1UdIVzzrfKonh
Pw4AdR3rWLyiD7houdrZROrOlAfaPnTb3pbvVSyOGJO4fBYqC1MseFA9CKSx9t+bXSELUb3L1XB1
phpnrbt1RZ/2N7QnKWoEZo3sr3qDw8Uz/r4pCxdOYSNc+wYCGJBe6HQgNPc7RCQjFMRfMFn7JwPa
Q0l0RCR+SZelF7ssW/tNwbkrm+/LT4npNI+hbAj9acQt2lX/xwZ08IK6MmQCG2kTg29fgU6lWkfd
fNuKfwJR9jcO3nHrkmZuMeJ5C7DyeXT3crn/Fh4EmBUTpFWwEbVf5fu7FtASuTub7iPUG/frMTOy
GxvonGPB+i2dUMAJ59CPWlEB4tvuVW+sORC+sPcM1UgiGA8//4wnkUh99f3rZ+jEA4qaJLctQ8CZ
W3lpg+FjIlLUAJFLnywV/ut52Z0/aFzM/7If6NG3aVCyHnITAMoJ1RtgaIbjXC9tMgQ7yFvU3EV1
svpmAvrcYFssyx7x3YhJvIOEZDc0/48Wxpf6rYmOYaUpSRRaN7jEaeRLymz6+KjoBqn3WibKJLw4
xnzX6C77Gm7Rqhh+cqZyLF5JNI2aG5pIjgSHZbJv3+73omweIoC2oCTZaXQL9JELpJFT8Sdfidz9
Txnrw85L4zhW922Lhl4Wy00L309doqbbyYaE64QaM5/iYGVE1yrNrj/debsYwEbNzMA8cAEDS1KD
B24xM8esl7m8rlxj36d2WWxGkgMswBdKw7I9S0uUEIVewEM3fuPMGvT4qmckzSkz5in6tkaY/Py7
Nu3De6C6uvLa7NYD5iTuOFqiDrbheNNCjlWuVCu3UnWcDwukbxnAdvvN141ZZCCh1/O9Ci6hrmBl
Aw9NOjeLEwXCthNpOjlDTfTT6lRTIwtCaoQMTdQzipJBDpfRKdRqUHM8h8i0NIoox7bvInx8CunI
zASbElKMUoA2UvKbZPN3GdD4sZOKHbtgO2UDSB+2dZ/aGZfCoAXurNRBq2vh98mEZeZE2XzMtRM8
mdF/+/DAOgpnjIAFUgKlopEaOjEm8QEGrdIr9eZNgrVgrLc+NxhjLjXzT1lv/crFp6aE+Odj33dv
ylnAijiQAP3hNo0oyZoyrfwisPbA1F9vUq+pqpGMybFejxfyFCYWjiM3B3dRsf10l6sHHxJOPbmS
cz98TD1+rwm3KrwlPk16RYqXaqazQ50ZO5UiYtONU1SKz8+dWWKirVDff0/UHCn/+V0uA/lo9Ygn
vb17yDgsNUKs6zo243Q2bDs74mpnYC8PINgkPWEzdvzp/WEeT1LwYUAwO576O+/3SY6FTztXCwkU
/KvLa+bSELC6UFf/7JkXHY5dTJbRVWQj7CVVxJIyz8TPNtebLxnyURk1MOdYKWUAnYfEw5jfvRQV
wQsYoMf4vnhAR5qSv5su3OogQemAKv/PgoCDtKWWKV8T38VKyh0MYwNvIUNXg/4LP6EoktIlFNJy
yrW9Sg6o9JDBbHChFC0boA+XRHK1nkyWNzrqT7p/YgZmSoYqOuBzQpw5KzATFg4Dij12E+hNC9Lx
Z4a8F5/hIvQtOPqmZXVSUSEn8YMmqxgORUtYs2H9ML1/ye2RxqpVViWcK8pOCXLKETD12itAI9Mi
Cwk7nBkHNi3AFXGP+coo9i7zTsrLfq/EctQXAlAQ3ODquhcSV9hxOTUAbNX9vRy8SjjJ7LTTKjSg
NF22iNVLTX9QbtY1qj6BbEJYFdFsEL/gDD9EcTq/UnNBANZgxHOgRji6bGgGHT74erVMv6jtieYY
28PzPsxX81jxF+j7Rb9sP+y6qH1NwtohIVJw2mnKaze47Js+Hc7ckZT485mrQwE7jgDasbuogFDG
6xan7u/7AV/Ac5iVXcK/mXonSBjugolIoz/T2vhcwJtcJcIQ6naTdXHXKSPsl0Pz+PkFS/vcI3Vv
xINMKfl9MmlC2JmBYtW5X0fc8g0cKomRm27AvJrFnMjESMhoyMSJFfs9Yxjpayo8NENh3rwzH2oC
6xsjfCzDWv2jTnHPIEqr0Q5T5xIGlgl/sITky88DoQ/m3cmHPyRifE+g5j0rULZw+Aic9E2IIUWr
QNZgOEh9ElyZYGRBTUOJxSDvrjORkQHfRj4BKaNvomjr92Lutf9G7hPpP6JNEbsbC3uCaZ9pske4
7EFeNqhLeKtLJcffYz/9yynvUay91HHoNRZ9CJjo6eAjKCkjMWOMoIInkic4zkQjgHbWbjyDoxcg
SxDAxj/QVZKNQiixYeKm+jDb1VaivGOpDD8Z23uP6Ku6B7LOsk82L5YU8UczzdHiO/pZVi/lu/uT
SWt+eeQvsA2YBAvftyHTOp/bxnIOXaNPM0h3cYnl3KHxDBx6tvGjQTWo3wiUSHpcisn97k+Zp4Up
0gqzcW+3ien8FRMfla4A4LKZ1l+xU9IbBcMY2AyO3W3BMy6qD6l3HHt+3QJVgt4uLY/EZHSwHFFI
Y13Nml31VUg7FOmHGmt0a8g+6zoVF6TXJHbh2niBJq2eDa3vp5uZGy6C+2c4jkHsUyEOufLgQb+u
zgg3/XyGqIUgdXt0lRl0vT0EfY06C+IglaZRoNYegs1E/2fKw/kVwTMGCq9MbRQQFrB8tYp9aaC/
Ixfd4KLeBfgJWhdjL/SO3qV7kOGpvSgErYvze3zi3880MMdGwIRq82fNbiZ9NF9z2TLCAix9kjAJ
qgIT+QDkpmPuGvWeIwF+vAN+IOfXMVI2zOOLRTrf7bGFMNFfUauzHAcel/W0t1hXZt9UN/tbqYPp
B6cOQkQfu2+XFPa3g2KHsr0WC3dcAC4wZXFAWPKvolnkP11vweXpPi8ySXkOWAWOo9WhqqGP5mIJ
cv1gcNJ+dX0lmX45YodV2kNwcVgPvuSsiF66ItWSiewjP9n67GK9LhRkv1JqI4Lr08Yjecf+Urs6
OaXsd+jCdfQxj1XIie2tIp59UChsVLTM8CemNJAtbJSZmpUlZjjmghZ1JBWhH9nVfR+Dm1uJWONU
F+Ji86zJWaqJgUvA+XJmjr5NMVotVcK8NWPQCtONm5eITR98nYV7fvP+BXNJSfDy3lWFmLSoZwUJ
+UdOhEg0L/IvmRr6vqA4eidAPMDzzwptgdfIC+/DGQqOyxTk0FgyrYR6EwoJI8oBRMEgzXc4oi8W
jznaYqKI0VXNJh+n6xKE5BBY9Db73ZwGq/UigM6sV2XyKKo0Le3UApq9aO7hTtmeZMTWFJuhexGl
V6hDBEd6He2eYrGbIRWRv+bRqh/747t/MOzl3wB7kDQtBbMJEYhUrCB3TJu7Mm1HhAp/3t1jR6Rj
FMrU98TaRYpFTgOsdD2gmSO3FsfDwmWUEpA0++905jAmnPqIxHGDCOsr4Qigy+/ouDt+foBMsXoo
vTu3zRvoSNef8F5OtMMtl6jwX3mppKC+/n1zWJTJAUf1jcE3Nr+dfOyWktEkJRPTHFseQbd0vepl
uGPVotf30tScJt5TFRZTQuHb18dBhpNSiQ5DtoKb5l6FCeprkT1p3JHrBxw1ckj9hZalmkzpZguu
5YHCYw07YtR8gHtIpk2+qdhB/yMXma55PfgpgiziabXwDzkqqLYv4JXupjUkpRa43jOtQEdVKqw4
AXR1YoNOiDwjDiyaLVc/X6ijALI4xsH+4lnxKGi6kpBh/fUv4uGtTV6/XQ5wcYSFBmarX1EbLvmB
7dd1zvwENZkf+bS63FqTMFN9LUmUHfpeR8DIWZJusk6GxLSrIE01kKEdditkRBb6IqPBgIGUS89n
zoZapIQvooVSf29VL+JphA5No3ohpZ5ZrGGbwVz7RES9owqclWi+LujPYknu+L4jWGp2NO05PSe6
ZF7Nehr5cbPGTKyaeY2qv3zVATyyCY3AiD8UF+O6fMwC2bOLcJ+8ED1oMAPlHlMr39oMAWdBP0cV
ocSn480XrvUF2Bq0R/4HsARWI1yS5Ag7YnwIwIWnDe8JLeX+4KatO6QfTcIbSE2Tq2pwd2h8WgAU
j55hIjWW6b06toeOjxFs4gFkORc3q8Z2iSt4hL+iFeo3UU0YH6gt//nMn1m0596SEmnt0tzZtQEf
5txs6KXv7FBThCU7do2zQFJDS9JcTCD9D1Vgu9snOfyps2nkaQ9UUEdLS7nCi1JRTDvOu00UEG2f
rcD4axGQuRA3bOxW/NlY0wlvqueBewau9NNTnbq3DQXIECWpgxxLjfr4S3ly/XIBi7JZfMUIy1kd
dXoAMYfwEosZC8tirGC+VwsAvZo0B39bcIMCPvNYWlJmWgjLgy/tVUzPb6YOn6VKy9AwgPrfNzzL
8DYu8ZKPHy2ax/d59Bs1erQnMAFfdcBbKWpguKEiprodR1smZr7v+BoQrrtsff2ct4JM9eGACTNk
kq/oU/n5N6gI6ZCDEG+02MUSJ8lqiRFJUpxqKDGV6DEx9unmh/jJxXPfcn3ig5safTP8F8TaYUUp
Oz0qFJcKf2jVyXVUm2A4CVe3BnX1u6gDq7toFyn/edXQYuhiQjMovInrdjPmTcL/CEsCL9kP37dn
C+uEowfY3iF1/3lJYMqf8CSwxVHZtgYY6M62cK5K25cHE8cUh6wAzzf69mjerUn8RnEhRsWUmGY1
iLcVz6JiHoEYjsReMjoEXXRJAjMvRKMQQeLsfOoFnDVuVZuaOvuJc3mT92gRwjxd+Eqo5tDZx8nt
g/BeEN9d3dvCTsrsqGWAKiT6MvrXYJFwjWfFEPRvlPhTRR6nPUbDBRcjmJ5EMWtH0I6qKsj34HR0
op3NcGiNGQRJAln+XoqRbGqAsUgzLyLxuBMIGvX2ZVQB1nYiEg7ZKL9OkUXYnccc4qCKtpBfzluM
qM+m9yGHHXXZvdPR8EcadpLdBW69ej5utWnEsY6PQMUHleWDjvYdEzy18xWv/Xg7O5/7F/KGVwHf
JZzGPq4frEsu2K7Gf1rCZq/O/yhwkcG13bVAx5tA9OkBxHoP2zsa+D3hZryqaFwhP3OsP/sDs1xo
NxuOYQQRLxNv6cYmkMclMlHb2Bmml7o6oegyr6m4k5muc7wcIJ0GWszEwTYpWgNLjQrv3p66I22l
8x7IUXKm1cedOAUddPYqOA10iLPoWBUJxhuX0O6hwfxqXde3EJaiQ6mcHFQnnBgXuVKbC4Ig3KcL
PhGezOHzbyolc/zbV5WFxJ8Sog2UQDWNimLUnFxMQJ92AGmRDsDOw+KYoYg6QfyIU8VjUDhLlAuv
MuGhvN/UbGqjxdtegLmU/iaYUyHn0/NKo+m+4EWvCoxLN1Gb3VzLkNQvf5KHevXx8vUnh9r895lz
OK6NnNQqShpbVPycGetgW2Fjbkcx7yOm8KY3c+cKjQjwrH3MexkLPCUpoSf+YIKI6V2vcNthq/x/
JOsGHud+XzOcKrjY9odzkkTYs9eEtkvFPlgx/gZv2hODfKIMCxUX8dUr6+xyEbOEx7EjH+4TD36O
cdk06glHQmk1hkYqzEBP/1l98FriNs4ZfxZY13gtFKRRU7CS8KXrsjt/2uKhokqzgv9YdG/uMiyC
daqTwXnFegErJxGxS+3RNeoHmZFvMZsCwPZ6tyqtUg7TkS7LxbxULq+6tmLgHLXshL5csPc0Fltv
ju6GJc97VrFgmpL00cJE/4svFbb0gWZHKMVSMjV7ZBhkRxod0bROFIxbd4/+iObYsmL5/f0xJ3Ep
3+1W3zxIAu6NyxBQhgvTuSKRmLvo0MUnXMDfBfCUTNl8ygv+nVo+WI3pfedP1x2k/2+zpVA5qwVC
AuygDYT05whplZ27+efB/cIZ9eb1F46k8MjuvRcz9CTXGAC3rRpbxr6bKocZ+dGkihvvsI9efSVh
H3RVvqgO82jhD/5I/Ex5GKyQ4hg1p5cUyNAUM0kMwMcQmpPvE2DVVjTFyT4uc7TJUdcN+KLaPGa7
oeLl8/A4OzB7C5bOisAQm9GxrU1eKbm3K8WQSj1dgw8JPHPqvszb8ertQ3TusjvACINfKesOMPVm
wK8S5/iKghRe271MswSywmyW04NRcWkqZ+VgzxBDxHl7QrSwcpOXnYHHKkUiwj7w7oRRUxT1M9/X
Yn+mbXJv+OAoFW64Vvz/kzymIbeqykfBS7kkan3I8lWCpJ7ccTL8Rf+37tYV1B+FRLvNk49rk3el
JxyIPMwmNIzsDz5gqxgvUdWAT1HhZsMPJ5YmIQHlU5p5/9BX0ANWs4tPO162A7dhuYXU0SJmXhB/
hYVmJK109MzGMsoqIiw8lW3JYJulK8q9vfc3Q2JCQyqg0KrgwoxDdSkdbty1gOF/KjosHHCyK63N
cHabimq3dwg63H6idGR29X8QtImNEXbSLNNT6AeH/kYKYEL52f1X6BcJ5OAYSW4J/z3SYghWgh0F
4sy+zx1HxfzQYbsVlG8U4cCPNNlQgMmIyBkkbKPdyBeqqozZKtV2gqI8enETexF4EVjqnGHO0anq
984Jd/6POR9fSkKC3rxtFm6C3ovSfFH/rievq+obnxs+RdysRhA1hchAOBSQJ0oRvUCszDudxWfr
NJ9ZzIqleBPb0oYuUJhQuHSGckOrg+bcb7VBr5qNdUtXztPx9qKrH427Px/UBFhgi7lZY/gmXYY1
WZUc05WDgE07WTrYodC9jlRHKJxyxY4Nj9HtfhVJCmcs+AHKBKDIllWzML2J9EUMLBPnaA6Ta56J
d9J+6aMl31v1X4CJnp62FxvfxILg+Z6r9Zyo0gF20wYOUYkXipCm+ktLK3fdpmvKEUyz+h0zxO8y
ttfdCHuDE+EXSY9agMc/Tj87KJV2X6pwZfEWMlsBxoL0d2UdibdJbpoF6k4QKiDJ9up7+fKo3oED
lgYVGmEKGAotAp1svadu2qK+rqceQC8PxoN2qq5FeA+C3QYNhjzc+ZtxqyZiR6zrLrBz4zdNIR42
NBqaafFE0hzoL0SWgfxHK0KwG3I+TFUg7uGXoe9fS0nm3da4WcoWa7YM4PpDMHvLoYo0X5heXW+F
uCRhTCYkV0GK6F0QMebG89dZ+9VkrCXzFS8DTbPf63rlS0/tVn7wZuZITy9eZ1bR63P3te9w60+i
mWyubHv3B4E8AOraVJC+hkyVNU576iJs/tFDTrd/iVPe+N5m0s0HLazCEKcnCao8YjQQZDXjH8HU
+jJGGKq3tY+Mg4KNmk+BT+B1lInWd6euEyCrIaJyBhMyblb1pvsP59DNTOPCEMwxovVC3D4kPWdA
63HwgBbh/wEfT16gyh4duBF1oaCSgjeTx6yzEmH7A9K94N1AZ1PULKz3ti9LN4sD9yvIJIRgGNr9
aCvlyUebmcFX4lGHL9zB/XBaoNIbRCFO8OHf9clO/sv8Dz07OdDGPfj+RqihjVTu1TgLGu4Ab747
WUCDAkdG0of+2ECv7kCVQf7HQuihEuPtIGA6DYIfPybN4T2XlHHWFZUIjEjg2PGqLWqUR6/oH7P7
EWsSP5xeRIiZ2CxJ63flL16YOz2Y3cV5jPb2PtDXG51q5DrUV8ix2yg1U2GULuXWug6nXV33hPbo
LuRfig5zx7xIWFIvSPf2Lftp8CdzJAUzk8i86pC+x00AUwW9ZjfdQMoKk5QDtDD6qRqwBnKZCHcI
gXrklNRIiY7YdIZGV55tTF+wyQhqHPRqfMWRNLaFZsXnagiPF/Tx3ZzgbGcAw0Ppdr/JuwpIGP1M
UbToIEC9Mm5OPiHxaOxo85xmCfNDrtiEXO96BDUm2v2B0OnfUDsmTz5f8kG6dj/vWd/3tvCwPDog
h4Z+9kaDWlbdXQSmB+WAz+hWVK9G91mgyo0rehh5cycBRfiqhakyDnS95badZpwVht/qNqwkY7H0
nmw8osaMRRzvxgfZvebKgkEQV+W1JiweDFJWhoj9FW4dtiR8KTMOgvY3/pvW+LET0+luX15PifOK
VNPllzi0zJQk7J/Cim0Qz+x2gYnR/BqvNb58EmnWKKojY/++pK3MVj7Qtl6l1NiowXQ+SCAnKRjC
BVRbNPMKNLP9D4XjtHyVUocZTzIk3OnhnVccyNiWGQIxhojDMf2PAW21mDe5DwUnft5oIev579eJ
SpxgnUnhK6ZdCUdZS+4lyWQz8xVGjk7O5cXls07ihLDJe948+NRQuUbiss/hAbWFMs6Fz96tWyk4
ySjmhNBBPmV4MGdtvjrMf0+xGSA0Z+heLBvTe9y9Y7OqjzkFpY/IGHMn7VRgXgWVSvwbrmKzkZ/E
lD7UnTmwHJq/ceD+d53QuP1923ysRsdSMvDoAzHi2fmsvpyznm4Vms/6oYZ7I9+7hfjj9ZeKp4ZJ
Zqzzcm+dEBAwhzJo28l8lg1inI3pBII4ztO07s07Va2KKA6RGJTh5VVwMC1k348Wk2+4ri9Y60HV
WMcelBeOU8WdSC1drwdQhezvKSn8b3k7YW7xzkRKHpRT8X2ZuYRdWWaoEfwqSeo/TaPGD5nqbv2S
GoS5eRYvCg49VNP0f4pVQXJR9EbyKJh+9SpLrecZE4cYRaXL/poVpK75Q9PfQUvCwo06lbo3KEKN
Vh54HfxSdeBvk/E/nSYGWWFJooUW5bKOSQK8VGx7fmrmrenAK6t9nUHBTlWuW3sUa+zbGdgsPy7m
k901NgtdRPa0BMDgrUePIAfURMt7OzztCmHKCD4sJ/jqlNTRxycPDbXmefYGF59Ee8hLTSBO7gac
SNGiXy4z650dLeiKmz3tGH61uOPoOfSQPKEuGJKSx/PsMh4aONZwqPcy8R3xGWrdFGZXFnZkm1hC
SNcCpRjq/0dPmt0Fn9f5LuW+88b1z1RN65dwbPES50qdz8JYtmxA3xcw8EG6xr1r+gAnoVOz+qQE
sAq24zf6gOudN5UXj7b0G98T/HwG2+N5LhPAoGNsBpynhvCClap7ARoDteJuBADEyfNRf/2+D2Ps
yLFtXOb9pfp2jNwOgwCCdHsOQ2w8Mae/agbBXGau1iDJkGomne9hbLp7EtAcdlF1w8nPbsaQ0v6t
T637v9UMnHwGPSzzvft6Sy8X2bofvakNABUgL51+Au3Vcd3AgAfrC3gYqRDuTJ4dwlTwESVZo4ZF
MrsCk6XHGwfYfUYZi1NK8pB7THkNI5gze0HS4/nYRDK/sPLvstDq+43JyEWOvsqdipf3F/UXZwRc
CB2gOf106BXApIbdJSSgVvuPN2MOULGSaK1aZelzHTE/zLmRMa+AT7ndluH+3tbL8clxG6cLge3v
F3qzNq9dyNM3Nh1bIsTdenuY8koyQAY/GUMtMM1eGooi69JCQRxWJQDD1Jqvy8hablEQtBEgFYnN
9kYgz+dhstU5DmAZFBtwujuor9dLmDat3frHX16GL/fJIhpVzXIyCObPbcUs1PyWMyjnAr4HBMw5
3vEaCdQvsghNfvQrGnPCftvvFFdlYJx+zocad7QS+ob7hX+on40mo2FIvhwhfoXUH3WZVqdSRYJw
5I4pFXilc8u1tSFCMHhBzHWn5esXlHJYSdKeaI24BjDBL8OTf1qB3fSfyIVfKAjtzyO4ZQ3b5fud
57KHdKs+Imd77syoS4WgzUl7QQQtG7okjVUT+3MB1Fuqvi1p2rljqzoT1+OAu4DuMHQJOaBBiGKn
JwCOwGZba4F2bP0sDa++IWICLbDaoX3i/V7KazeWAxPYLfXqj6B54FGBYUKnrTXK1oa8AB8R4nbw
EvzbHStD/d5L0tjG4NYR2HgjN1W0moSmk4Tld/2Ob7z7GeVV8KFm3lzym4tNL0cYUcPRI3q7eAkH
FYAwl6N+6JIitUjsL083J5yGk8ta34/aDcOcCXayVafDlf5P6OQsaWrj0mP6NmLYF5OknKCpJOf9
AuixstS8KecmvH1AzKk1n0tf3Mn+SdbMRT2qAUWB1Yc8vwepJkJE+2ad8Kdebi9i1PDOULF6ZkN1
r9sH4jkgjhgRuMRMzXLgFCWFBNgDDCaz4tnMZ9G019KHC5OZf1zyVucITwTkiP3oBlfjmCXi408S
tci7pbqkOswDfG78wHnmuwX9nSCkoXPc3imnV6YLefPK0NtgvO+L4pFWKVY3pBh13pq5w0RFGIkD
xt6K5bXQ3SIwa7UYZT2iJRkEqu9HDdEoMwwG9jhiZvZ5q2Ee4QlKEiTURQ5dTyMiuxCXChXTe4Vb
XUcU3qpgPIRZ8g3NFnWq9+RaNn/o+3Dlg6ZdYGpvAl6zL/vIz1v6m4pS88IsXb2VBTHaClBboWNO
XR72AtzFwSOqBYeN2lEjon4H5K2Y5+e+C3KdvLBvI44O1sCnKouEDvuSIAq8FBBUHemfaq89tBXG
pxx81P3V+yHvNY8fxSN4zX/FSwoB7PRj58yIWw5r17/17bpdQCx4EWdNYuKT8/JGNkNF38yRzBk8
lO8VQwx2cj9jPL+T9Q8eV6oJMwG/+3ft0rCaYsrs0aILQU4CZ5Y7/lC4gYoG64HvjmzTC3frvQI2
LKpotHDxLFxE01WOeHP+omivoPbSef/tmZmG0UTHazGlLHrSEUxwSjETzgUYNh/QkvpauOS69kGi
LZe+8nKzn1wFEFoS02MXksYDB1620JnOT9jF03BK1FzlyuVtNE39RXmuuX4U988qdedBhJ7m5inB
34EXR1rksdYGRuxCGsGOkfxDZsNvwtisV8zxm0WS9mlwRXNLdQH3/YKSDrj/ANi+IPBYoW+k1LdA
BaVOyC/XDWIQfaDLTaJrWplZf3llDAFLYwvVk/VUrRC9VvA4wc9/bTWnrRgmacL7XpTkNw/gJ7aL
tEYDxRyX6mZplby5cyPRmNlTzg5Mg9dKqwP0LvGkUlVyoqW+txVCVD6oruP/qICLfOIu/+ATqRdJ
3vXWpks41GFs8qTDJTA8hy25HplvyqncbAGsz6zge1MVlLMTxAE/LgWli8y1no3SAI5rKEaKQyiE
8RclepvC0sUkWI36HTk0K77VCaWwABPLoN74hRCIKvlpuFlxpumbpvrvxzzp1tUyCGuAiabC8orF
hHrVOkg2PnSdAL7K76i8BlyIEPYh8nuc9FTLhxSYztikkujbRFd03opDPD9R0GwHERk1rcT+P2TX
Of2UUCi+bjmEUvGpD46A/vdJe2mqgaeINl+KqJP69hZqse5EYAPugDy26jWaAXKaBZ85psJSWuJK
aoWSzJs0x54cbrQ/AJrnwfONDSHSB2sp628dlXm6fu0tWbIijEtvO/QwuUB/eQQTxJ9ztJPdfCJh
uNPgqgSRME5hFW1jhq7kFAssoVSABRPA7VlYNJiGJtowroz6tdPDgErMuV1/6gQBGhUy3Fwj8Nlq
ARHUnkfvivmXYdQQsLyQHOfoC3UeNykI/GMWybbpHF7ZUT96IP+0QXh0RQXLSnK9r8JeG0oO/vC1
98iwd0yPTS6GC+3AK8oM+eOsKTQfA+jEoONkyau5mn6/lTTRJdR3+5bSam2iPnf9vb8Yp/63GSLc
F6xSdVW8Tp2Z4F4s2RTFjXBiOn38Ddao8DJWEFFXBaMmPDdfQFmGPqZMPfe60QpuOutlfQNHJNAZ
mrX6rdNwIP3ahyoGob9MUywTmun5wxfn784XU87uv77KuaC+0Wogfm1NIMHL8mcllJL2c7kl78TD
rmhIxp8iMI/Lkkonk9Pd49x0oAdSFXEIxI/6wSjgzaSKUMj4lD3goPfZVilgpiKL23LNCQuEm9U6
+Hf01bA3Y5c8yVNplZjITBw9PB/kdLgzXQQk09zc7KaoYgcsLFSl9athNDGv+iFPpDMf2qTTVEc4
Y5ufV1TK1qsKDuR+1uVu4BxLP4fDH/kRjyVk4CIiDyoEfwhEBJvtLY1hN2b1VnKyYiOdq1BN4bhr
0b61d5HErGMZE2tKpuLO8bGQrBWvqfxfNVv0WZsHDkvxe25AnWPbKWBpxLxHKjgAMbIFyr6QFTNR
vG9Ve+JMJFvma31opG4Hcw/kBwvnSMfB3lPZHG2y6sb8TII15HpJAgZo4Fac7woAyYzjvVtB8zgH
DtJVwW4hG/ZOX7KdO9DhzBMFJNK/f/VcLjra6XYYbqIBCP8HMTeyiIcC+p5Qm5HjTH03W5Rj1qOF
BCdiFwcTm+4GW/cLoUL9GWlek6YjTZLnAd9Ve9Qk37JZ2vlw2rRo2L44vUSwGAtsnXE0Nk9tGwLG
Fvx9ZiQ2uoV7C7CbpMq4f8/NOMHGvWpCHSIDRUeo0QOgzEKSoGQ4IpQ146I210hnRnyNwL2NMzjR
FZ/HcYsqm5UBmbAb3M/Guqfn7efgmHO6tFUfXLZCZQLeQsnaGwOLNOl1ByhDe7NeEXc/pn22VGv0
OkS2U0+qwKRmtxuMnPyzjLAdtFUPBvjJvbHv1WshcXDxCan0xroR0a1HyZxOi/wQ/db+28iIWq63
PqVlf/4inwsvhMOmMpEj/EEhxFVrCDeQUPwnciz9LijdGoG1nG2tZ4c4xlopmEQ48a7dQCtC2TVE
qNvpKmCBaiMYBxgAf34C0cFbhZ4+hQVhhsfjxwXDKOUnkkEoyKT034EwpV/0oGgzP14ia7LfA6c/
5pDFY8ZrhPAcWeMhUCT+2ismO1M5UWvvs/WlPzfaA62Exw4fyxVsyRrb8wMUKpi0Wba/4z+nulCw
oAZMF2Xi9MiYkAgCDfycmRClBMGaaEKUWeUWJqfqffBDRUgzeywNI3PuZQkv87d7EPEhlQWT+bI3
9Va2JSpvJhFtTv5I3YiqIIxlISEqpf6zcsOYoyap5iYYV1V1kDbu46OAkHx7T+TWACB8gRTVQ3vH
xnRX0tZ47gRIE+LiEnxX5Zacq0WLJQ6QgMKI9w+52x4aCRLRLHVE35x0AeXS6ZJ0w+aIIB4sfxCu
opBT/SzIM8UbAjijp6hc9UwalsaiR5nBy5emYDEqG5NQrYGJ6s2lpiFOY7DOqIvyrTDKPLEdpsFv
pqhy9oqf/d1MHSMFI87ajGcbe1UFXAHAgGIYoPh9rASje71nz/Z//CgPJQlCngG1yQr9epRIjbWe
JFOaEelE/XbaUpopDOtA8jgMZwJo2SA/xooyTuYZYtiOqAi/ItzQSCW9cAd6rw51eU2x0J6zSxMy
TlC3paVju2tYEczR4RutZ2EDfiXnPhA60Ibgr5FRL6o00++STRjrGfmbX78zjgmaiqeH2HeeROcu
CTngauIMnGdCtJmjZ/aOS8Cx+aGdD4CIUrd6krMd/nJlmdmXZTifGk4MlDM24j1bPkYEksIFeBz6
M0dj9iAdnvTTtNLEJGheNEU+JeT+13Y8SYDov2lhBQ10rQfxjHqHJ7MaFZ3SQp7yWrKCSLWch/TK
YgagrCbAoGQi+JswYrk4WaA6iKSRITI5vel5rpMqfYtSWp7HGqkX3Ri1KOyk1mrmAukMTISfUZwV
2BhnQdB9cLOwkMMUwkX0e93G3Hs4fZPzsfFEdPAzefOOxjT+4pS3TYtERk5T49vAutxRWD+9ePoS
+fIBUawiXtB0ogNfWDsM/ZOfDEc9wAD9keAywdSBVU1Pb8dnfmK0yIeuVQ4CuSpmNpPjtAuckmrR
Z7S/1Ojfnnbqj02C4z00ub2L9nO7ZzLed/aZhBTfXaO6IpSgN3e9jxos0VALDpbqNQ4vkCwXqlsZ
AoVzNDMCimskBqPr0F5IPVNwtqQCyDsWsukR0k9Yl5r0syfIiaWrSGebI6qJNrtTbaMVsSk2BD1h
AOukImoi9//XzGJbVUvl6SiCh0+XiDXiv6lMAQz0RqB7g8ERtnP1n3I8jCO1I3hdNK/EezmtWnpn
3ZAbV6EEJscC6qwO1BWezF45eDJ+LcUE3xLHjKFKQiZA9zxVawhw/F9/h6sDWAgVwvlzMR4H8E2b
MO/KiSsaSqaGkNn0cc1BnKzjB/6lwPBb3eOaH03WV9ZrChksn7+Wi395t2rbBXp/3Sr8+wlhtusn
L02wCiz7KwywzMB7wPwY2KAuh2OIbg2eDcttMdBPYDhHTR8lqeHABvk2dKevpQfZxednshEk1Zvk
/rxMZVmfOaOSZpE51k2VkSOg/YemsLnxrZH7X+0WEFtmTlTNB5e2vGjtpnQ1vuCsL+tiqncdsLZi
EaZGFtsLCCkWRggWaat/0ZdsNpAz20FNa8eKpqxJ//A6qT5k0KdCFSMQZOZ6kozieJYL8Jm7P0dP
cjHCCDQj5ajuCRqQeNWGoJ7xDUEhQG3q/iE5RmLOwByYCGEN75xOClozHpZtpMEJ0TEMurJouAu9
fC+ifKRHRpCCSrYFyJkjh59w0UagTFGo5jecEmhYpn399C4gXPN3S7kLdcl6JGgRwnz003Le5C9y
9rij2gI66extDyjW/ec/M+j7kuafcJGMeTcWh4btmcmApxaGW8HE42l51B6Qm70fD2VVcRtOrqx0
waAL7f39YPdY3qIV9WWWZiHz7pFX5+VH0zeE9+Lz0rjHTALcuGW3m0FYpB3nwz3xFv8PN1ODBIOn
kFVxxLLXDOzaY+Asor9wGvG+0wqtyqaYPBD0R+BP9I+03xuc2VqUlHU/iWfUapt1Ghoo85zoRZVy
zcTUq45nQFcRJcMi7FH1LoJdPM6dww73ky4HdwoAq2vqjcdnig/jS+cxvpP7tHBBjbniayhIjqKb
EvmfAAnvYpXMsF955VfBs43WWh/oIifZ6z32vIyumAnaf8XcEy9Qp8OvhazCFjyKwQYtmK6Bx4yk
POaBtSBv+9aU4BrN5ThBrDKgzo4SBpM+27mNX4VQC6OnE/F7k58pg0M24CERZkDd5lmiUYJfCTxQ
Nqj1226Ow4KmvmcfyIfgFnMlVBrG+xANpbnhBjYF4p3gAOnIuEE1uwplPf9tuVUx/W/kOQ+/znrs
oEuS6I/hBIYq3s1L7dPd8zJVEPzmp3ZOpvZq/JdOULH9uebdVcCP1XQ5l0yZjYccpfeR1p92zPhr
L48g5MMFqfryugPIcxSwV0030TasgmgJytBzbDRliHM0uA0A9xHySlpGlAMf300RMdUsJSsGYS6f
9zEDuo4sveIYQHs1fhMmJkNt/LimeL+bB9kFObjQf4OCbH2Ni1jTR32sEiidoaOAJInlXxNvWwpm
R8T8CuYnTMm1ddcjBh5TrRtrp7TAPrf/6KYs3cxcgrTQzzkrK30hDQdJ3SfmETm7XUID+2Z5OeBX
vIHhHDYjqdKSlrtsA/MhQUbch/MhCpx6d6AvkdUKj5zzv88j3Tu6bE/hEMAXhxMnqV/D+lTc5iuf
eU5vC30CBqWWBvuHZachK07sRjWx72nnnL/I4ud0VD/jJWPo4nJjJ+Es2S+K3XNwhez1ax/acTgH
sXb1DNs/uLlBKE1H0ujHQZXmlVmIByd2+fagncYX8nFwZqJGWRSVne9Pq9TmAwUNf3etuIN4OIdy
tCjJVQayBZH8mf9aHKLB8Mk7LAX2AG+SQuPCM8dcjo7AagETcZl5JIwltYCOOGABL2x44m0hTuru
CI03i7xGQZCMSbYD/VO0oGmnXSx8M5U2zZJEdnNlt2VBVuQp1KKuYZKWiEXZyz90B/KSm9Pjr/ff
EwmgsdoteKV4OKFZJrW44ODk+ejGVheOd2o/NW8RLjSK7fzcgGfJxtTXWMCWQQqTMeEg65MdsFEP
LS1HlyLROesoHYmEtguaWEtbbKFHQka3oTi9Ps8Z3rXzrdgBC3VOU5cCwO/JiIodUcgQLxx/m0/k
U6Ht5JS+1MQ182qQPap0/NFv/+9V6mioPvr5aKRq+Y+LIYfCWXL4MPGfh0cIqF/yC/R4PMy7wq5g
01YJQsLGIUrc5qRG5hTmO5ca3RGxN03TiWhZZd/ZboJLsoJfJjkuAi7Sw8VRAbsb1F0dIEnnqqKX
0L0cdjRwXQXr9NBaCB2++70yOe3O1vsQTKCiUEWCA1YEXdpTTmsJ8BtTM2u1cN4yx2GKdMBE/2+T
aKC3zc+r5xXzs0LCU0tyNMxKELEZ0KSS437r+mHgwTzRWauu+9Yxhh81pvqaCg88b4/pQEWYBZUt
koonQBGF7SE8aGb/MvLW1DRutHw2PXxu8wf3JS/pbrgcVfyIOJmU7HUyBauOWYAqF0WDkkCh5CR7
FnPMK4CKtydCHBydvUZASN6XmIvWKc+wMxQ/dmRQNLMDeHIdxWFUnzSWlgKIE41gYyMbCGvBHhbw
9ihTzqZS/9zmfLiTV11meBmJflFxrkqDfa56np4JUprwUpmemFc4HYLSKZJCgSr9H20Bktk77T/g
EUbHA2/YdtW5drZ/vrQmLLdWUOqoemtGRQw3RedlN2ndcAdeaKJdNK8hmVmR2vdVPxky4UNwW6jw
a0hjSMxy5pdlEzZA5v7lW8AqWWm3KNcTeiiWysHfow7VzYyVfhDBDhLwU0V/mleS+Z1aUlb7DTO/
OI8yssrkr9buFvtYv9GDigikFWQ6+sKBeiSM5QPMMLkmdMqird6bBYibezflqZy96G+9puMQx3kz
8rKn1b5EMoOicoTTDncYzRWK6hSGwk2suw5ptpM8JsujTsf9O7GLSjSky1p1Sy3qzijY+efaWvJR
Ewv52XO7cWi8c9/979UkCihX9/WIG9CNWWbOttEGpr6RQKzyQlQjTBjLaJ3Yuw9/CmgJyR0UkKiM
wZWtZwGk+u5q5RpkjHLJDJHl6oUK9iFM+kdHznhpfxp0dWYdzZeYZU6k+96m9Nh4ONkoxFO2CcD5
iLFAD/nXH8jESE3eR6fnjjFRASAHz8Mv/wcXaOmnPxYA3KQhubnf8TnPhR/dy5tzjecgbod7AZuo
zWuPkvCmQ7tv9k4XAZhKLfF6tINaPNTMqwbpkcaDWT6Pr86sFh75HAkAO+CZMqxl06PnA3SW/qwX
VFpIV1A3H12o2KWQAAdmTWOHcde1aqJsxUBaMPraF+bpzEXJQYncK1P5NXNwu43tbww0pOIvXaNi
ZL3I7z0H3eAkylD2yM1gSH2E5kVMUI9Y7qpztRwc1sHSCOSj4OUzkaBHuZOZfnFZw0H/y9Q5fWFK
KdqEAfQhV6LoQq3IefwUXyGPBFUC2sSvfd5pOI+13Wmz79ZQLvq7e+nMQQfoBzu5zikCTbWMp2An
uA6tcu0zueJyF8YgQHBWfKt6QvuWjmfzRu747yxDC/4Yd7avMWLHDq60qB9OZ8hG9surGh/HfPBc
7RVyrExYn1GSh6QdV4uR//NawTp/zhMx9FyI1B46iehureS29o/sbRETH6F+TA+Yk7PjCWnkrD/N
yIcL+7xFDUtOFgty2YYwfpy488vbXVEqXPHNPpMzYGlp8Q4IPYM7DaqYzgpVLFBlhz89YTTe8iKf
0MkYOVinPR8buPCYnKQf6ome/qiDoVDFXl7Y5RTmkF3WQNXfeTvr7kA/Rj7obMJuxRuRqprOiXfC
a6JWiqkkDNMJY/q4f4xUQYkPBQKiU0BW0OpgcXDPEYSKI5l4zhlkq1oHfZVWdthKRgwZAmHgxmjf
X2Bpaq3SMYKXt7rMn2f1my270dUS39IMz6mtVf+RuljVEa4wJDT9EcusRZJJdjkfYVwoFqVDOdhD
aDnmupVesV4/BPbxGhQiYQ9ObLK2kl3pyvUIImn6wul20oQnA8I2/1/rkormJ3mzB9oUyaY+Iq71
/tXvVt7kPQbL6VrYelEjztZG1Oj5KRZfRJPRcOIcLkmASGWh4zbnZiXV7SuztMe6ku6cvr0Fagh3
0OSRvgnlHiezvG3JK/bsiqtEpcYHgcmcRVWR/cGvwwiNR739V342zrht1dZ280LsHn9ko5yHXLjG
OQ7Hq96XZ6tcRb8LD53cdIXmT6tq+/Td3yQLFY7mS1q1hoNqELZo1tvfswJFv5VgE/LIYWHRe4rO
eWrnw+wSdm6THoltgbWZByJFqhM4PJ6qkHXco668fx8GXUsyXXjOvth7/VmzaYFDRI+oPa+9eVgw
wArAGk3NmPejUe10mH+qwW7kmZULLJ0b2A9gkvUXW9x75Wvss1jdDFkgd16OoNyOMUHs7QehPbw9
VuoQ7+ZIbqU6e2TmEh6H8qJwWjN/q/CXgXtqK8DWNHH1KyR9ccjAMWngQr5Xkv+qXAoezjmJ5SZN
cMDlXtfsoZGWpMyF7bPborICcdvLk0K7AgyKK0jW638R4r2kogj/7n49cAA8WDoBJ5v734owWQIC
RVPnvq9xm98JCkMmlTV0rXI56NuSU38LVRYyehYSzw/AXDDCzTrM1JUv2k0QCfqUHEMDhSMcqm50
xwXvK8lyZYjLS1LLTSxlZU1XGHvMl9n5RR7dnBaerCx9bWSYM7yJ/6Mc91o8OIc+/MHt3YyqFZ50
3A1DVjv6ry/ZSfdfvMPDujTIPSVla0nONDQsXS+LjtUZPrh/FvYegWf45t8bQiC871a98bWNl/pR
XeNMzxGIZRvmjSCIOrS/RJlNVcAdCeEejkf+RPiteDKwBETM+YNIrJHpd32iQ4bEMrIi2ygIBcXG
PrShvYvaV7so5jW9BspqaBmn+zCc3ZN37SZHHcpMtroWhU0fceKkezL8ABJmzy4+QX53aAhkKnyY
RtwsFfNzkXw3Wo2bps7AhQIgPbtcz0JjQ/tQY6kO+WeSiF03lieohdER3Z5nY94iR6ycERNNWCtb
beKz/UWcqYjYNsPa5dX4Q5ClY7AqvAULvbc/GsjOXfiECWnWS1XpezNdZ2jj2kMnD6C5lNkOi8sh
H5MNW/C/Dud8r2/Z5q2/j2grfz5FN5JkW/FRYnvZdLf+L9x7Og+IesbXQ4y4vM2JWrJ/Ey1s8oR1
iNKKB8dalfUXiehYLpjadtIMvrot+wBuHfE8KybPlxxgihUdpxnuDSaKuijLM+av+hyznB2/S3h0
KGix7l6Sws2ATuBO2AzNUzhxuqzjBziPuDAtIKnaB6g3+2ccOzS4fdElJo3gU0fQNy/gQ38/jpoD
4i1vv9FyNjt1jBcW0Gv+aFw0pPBNaKbB5VfSVmplzOT/gIeRg8VVGIfv5pt11raNVjol/a9IxF3O
nWp1bcWwFpBbnEPgxVtNmia1y9iefnlg+z4OwftYWYB+51mdqcsQje6EexMBaOgBkHlqJUa7Gcfs
ShAWQ+uIP2zxVwuUrexYFw1EHG7sGtr4pCzxZB5NePowOBv6ITIF281mHk91HR+5PYP0mV/6MI0/
59q4jxjbhi1kUHUNOKbW7VCwxktW52fMWfp7TP/NeOH/mnhWsOBVXgsvLnRP08tCPla9/IXAAUcz
GTqBFWxOQcbSgl+5BWylwuBpva8E1GK+0tmst9bWe0jDriTyWXpVoNORs+a5QoEK+oTyNBkMryJJ
JHusqenbM4ahwHvfwgSgX11MoC5F5IiBAnBf4ocBiEPfTHzlAMZZa02BKPeQH+IL/hnslN2bEOms
dY4ZfBBVPehKfnfp8P68xK+54x4PeYKr/hxTXzvloYjnOhhtXJlBAAdMN+xJVncv34BViFpJalWj
oswPlZ1fDMmvhw2mYro5wDMGLIFupz+lZHZO302aMTa4XX0NkESlJ3VD1E/sUXvm9ejpzG9gIFB7
Id5WRUyiLpcMeJzMk8YD2mRIIzTVZ6kPZ63ksnQo6PriZwsSwVAF+QpCJFypOXlDhIy9+q42uXRq
5ZmixYbp20wqQeV0OPohmFfF4dwrCtGpUExLmt7ly31i6ZtxayiXg5K6eqxGJstOLAqeaJHkOaio
aqgV7Cv7+ibmsj2Bp57i/+jYA8hWwz1AzJQhj9otWYYIxVj/vz66y99wAzMSTcdRhUSaMQ2obviP
kuFGoOvUIRaJqtQMhxxCoOyqe/SKLhLL6qKQnw77Wcevr82tlVGPpQo/4YE6VBuqiCPLps8hTsgS
ogI1CWSU+Dt7AgwAthYGrlYk3Ns9UnSsZI/paLp/DmAmJeCbsPAdUArC6NuqWzerhe1zRVroEznR
v2g78jTbNXIcMUv+/01HQIy7bJVsc7EiR5cZtRoLXE7pNOra/jU/TeJAd8NQkhmX6t82bBuXG+ai
Uh6EMpSSd2RsyiHyVWRr0EcQMj2YLaYvyUvAyve3SGZGB4a6AoDtiJCwl9H7T/ilFVFwpcIugE2A
d4af5GNkYu4avG1SqMoNC05hwcGUBP8DQ5phs15i6gAtg0iy9zvlkFlkNJszn7yfNgA5OMzIMl70
juFTFSRJT7P242KjBuTgOQj/kWP8UGoWWj+5GWWeaEvsBo/7bGBSl3CcOrKWss1PTjpT5hNZt2YC
ty7ctRF8y75Pbot4KjHtvZ92ZNtszVLuuR56kArYPmzGEVV4kcPqmz/+m3SNG0FXThL3dNUQI0Rt
EGx7L3ifeQLRVUakEpLoYFg/6EKJfdsqoaZUrZ8RuTQVRYosdPmCx5m8spzh9oDAWnDZ7X8c12Hq
H6jNYlKTrr9vqEwcFWp9uDhw/oe/+QW5xEzC2pY+FODcf5DT9mRLVtYzY/9ym8HmVYSKpRjOUl8P
0nmtUmuSXRwm9xQB/fFfq0cpEC500qdFr49cu4QlvetguswsJk6YJseFXGbX+9verPXuhZ/CK8bz
i/6MENIdKkpL5Hp87DoTiVU++7OesF3RWy2xwdK4rC6DPebwik9i22N6Vw94SDzzdUlb7ohOnWxF
UGN8PlH+tP36LS9zBwb6FEZbKZjy9owifwgRsroWsHbGi2eRIxhiI5dvO9x7Zuu35nK7syeD9PD5
C1ANqCYIdvrj41WLrpyD53hBBQIzJFCB4BsmvPz3ialEP/RCcUG7QECAAuWU6TA5jgA8MwF0lDHw
u5rz+yYwS21DKj93jPIF643mpzd59432Db7or8vG71duLZ8Q5JOCy9aCAPv0BSS9zvhigQ+ovlO9
3N8QTN3rPms/KsA0E7xkrgg9b/OvojxZLIEg8kgkY/3RyHGaap35kGbz3ofgwMIpIvzX98GN/xKM
TUXdI6nxXWr47RHet6bSoE9XPS8y7AZHQqkfXiagL25fHvOh12MNeHghrMZdRO3hj2w1ypuas5Ge
hGUgx6sU9XDXNQDW/4JIXziN6pknwAaH0yzjzepK2JVK+kuQ8uemdxrctPuihRjBSPGP7sbel3IX
urlu20ZNywiWv3B9StLUXqkHKtIFUMAPBdQOdrgz6Hbwqm85F6uLfj5FNHlih4G/P2GuHHWKHQrH
AsncufQ5seZAU/fV/5VvPDf3ccUaBlITnVKU4AFTC3J2l8i7u/Uqch5mUEWdT9uVBGS86vPDu1Sd
Rj12PeQ3AltaSI7PQ1y87L5MRMFILb0Yi1yXmr5E3FMmWHeq35ra+m6IK/fXPBlwWw2bi7W/L/yu
U3k/BLG8mQnd3bhuXcUOHvIeqBfeREx7DohwrAkbVjg/kiQWxFZbbvYsOSIgnJ67kBxLzNZnebpa
Cfoi81LzTnO65ZfZobySOkQYY9bNW1z2e8qW9AE3pqbilAiM3trvqUol0lJMD6mlVQ5yPILz/01V
tL/nMtk2NXliprqmccB6T/lZDKVJWtl7T+7Uz0B4WHhWEo2snjAR51I3lISP0YxZ4kDoOAey4AJY
5BR1Kqf1nIJYGNQw1Dr/Rsj5KoHVhoq9lPMQW7KBGZaOFjeo50Q7rIpSCgK34KiF1Tid77pK433p
uZ5LBKRtlVxhKKkA/zpJoge5+PlQ0A76ALUJGldKJa8pmNcZ8Cp1OGi9sSCjwmx9i7scRCzlUM8v
wGPMTMhyjOEIDlMTSNT42aSl5jiIfiVCpKpum6Q0skNFqN8Dl4yHBuBOLvcQlCQKJjYoMZFswE1w
5swhLCIHuO4dXlJBjSlNviORnQGlZxKEyphicGHUiOySavJHid5cZPnLBwuJW02C5zgj6DxCUErE
Bjdmdm+th4m0p0gyoN56ABhwmkql04bqmpmZsFFU1WbM/dWG6TyslKQ5PFt1TZe92PKfbULwwHuS
PyA9lKmfPkS+ZNq17YPgNBaxz7YnWQdFtzilb2ybmS796veFaw2JCrMDEffI/0hlTOyx18ZqEluv
kz8JBo1Urs15Ub2qbTT22z6Wf/vCyh9LiPYRIUOWovCnJA3tSg6PzIs62BVdTVguE0c1TrkGAoID
YffsoTbJuuXNYdVIysfdN/7WQBIh2ZDcpm9Llo0Kp4uaxv944Mg0fyBT30aNOiP/UGSlKJ4y0C8h
LXyc1Xf+281rGrKTZhDjYcO8d+5z3atCga9qddmd09oLAih8BxS0sSwEzb0wiDy2j7Vvi7IO7bFs
LA88dzGnXRMF0tnNxJ5L71CZY50csaHPnv9mDGmMFPy3P07+/NcsInWCcO8cKAv6Y3Y0e3ddddwP
iHIX54BgCwBPKvoaZqyKssI9FWT4XLGWZfYJddGw/gT82HL0cDFQN9izp/wP9DYUG9Bby8diFjFi
nSXouri2WRBuqu7UDzOiEoyqcHNo+pi9TcOAOHuCuf1Wixb+yX6HyLKcfFbAXIDuqqhmGoYuHpfi
nIkV1Dh/sWPnsJJzZeICH9rPw7ai969OrLV+sNUxTsNZWfzw6BqRvrBgn5OhDf3QXhOU3vtlShel
4J1vvSxHvEN/BoYSCyn9dZfeWvCNvtJlYPEFlIVNrXYE2Z+ab669IH1eqfanjBL3Sox8FobqXO1x
rpV2ZEGT9I0qcqy8APbIGitS8wfC6QliY3aPl9rwNtzgMi+CnTjFPER4TwIWN0auhHRWSrlgFeeM
lbFCcSiylVYnLwRBaJFJ/Dpkw9pB9uO3HCuoarCelP5h16fFICBB2r6Q7LxNFO6c5I1y0uaO98Hp
dowlFRJjG2UGyvn3cUggXY+1C5/XuuSzNHGbT41Ps3ExMjyWsNhNyfJX2C1hn6VbSzQoLcIIOgVk
lVlE1is3+Z50/oglxExudhmoTwkO5W8A+9vfbYM1m4vxw6ngzxBxWnSfP14KKgcabcFbxrY3iwQN
EAKSRo8XN6y7ZL6w+w2KncijsUjgpMmpGYblacqUE8ubJyeEgLFwpKLLofMWZNecKaGOK7Dr+/pj
0+Fe8c206Pu425gfIMusWQa+I8BtMFZ1g5KKjuyHymwP+l/mGqD1lBa0tGYcmfpeX+xKZkux12Ji
7YL/7gJkeBVU/7GsWhUlFIoQLR4QHQB2OY4nyzz+K3fdUf3Wi/Skpugwe7tPNPWSrIEn57Yv24iC
3+Q6nXVsjcRoW1KfBg5UfiN8kWsCFxhxRNKQs67w/YM1IZx9bUIOhYObkQ9KWjE4GMfcL22C+Wrl
hX8trIFcurlFNmSwH8TerjDmhlpfFabK3SrW0H0W2ge32gK6pEdNYhWAcwy4pa11EuowPTpvG7vk
z3NSPOeh5xEy5BhL3UVRQs5EzMZChd+TAarPXTCB58eItVxHIaO2SsSPqSb9MtB5B/ypElivBrqW
Q248NLN/GSC4Q+tgSwE3JFUzbXwbeNsvu1mfrdXXE/kuFCMSZygwk3drA5Gyyh1zna/fgoimPAJX
QoQ6L7xkMfniOWbRNoe4xqKP0+XcAyum6dBwCSxquYGN4wphecxK1mKEsqGKU0HhGmusV/cwRckK
YJfjcFJ+veaCR6ixkZbQ7RLRo1rpcAuooqul7NKRwqfrYOPgdekVP1/89BruKLHH3tcAtol5jca/
zHk0MBOEJfSAr7Z69ShFSSDbbDBuicHaLmlT1YkL/PwoddhgeQznQhUUh6gDSaKFO1dNPr3ZokCe
jcyJ1I5pyfVpFJ+LqD/o28HjYVwCo/rzY/fzKI898dH+4urZDTk+dPUSixslXElPrrOj8H17m6Id
0tvww1fy3T6p0FjX61BNLB4YEXUrJOBhYNfKqkVs0osHDKliRuWWtBte0n0QKgMJ8rPkEH4kmNfJ
VriiN/+odSAouaF5DeT3dRFb4Frr1zVbsAnOg0Yl5TLqqPFxq0nEw4nPDdpRnndUjC9WRZbwkMsP
JmysB2jZdELmezXfWrcOOVxnHoCl2WiLHIk5zN/xPu3XxrRkXPMTA2JhHSamPAJjU28EoFo+Qpvz
sosh51x8uu9/Y6EgEuNnHyQZ2cw3xsvXN57wgXq2PF/JwdpT10aLZoOIBEAYlcbmqkB0CJg15fUb
GbOAPCFi/rMHKBvE9/DNmR8q/ZQzgAgW/S92G5pmrJUY1k03FVAiaOnoB8RNajQ5HO3CVIys8iMw
B8nFxBKn7LMi+/4mRIkaOxaN5M4aLXBYtoc/OBBUnfwTuSIY0LCHmE+vjayPkf9Nwr+65TrCRUdk
OQc1uChu2SG6DfCrOCpjPzIwc36p1Ap/hedFtX/gVHRLg2EuXHUWs9IE9z5N+qCRInlpe7o1akFi
/cjaSF2AmRMiECXEin8sC7VS8wHJ6Kmp4wCUdUMIpaAMNLzvyQM/Wrwstvnh8QtUqb3IkEH8iMYf
KDIDtDcOqXzZBoli1/o6SNENJ8L/9v4JfyFkP0rxVhaJbj1mB8K/o1yxfU+3vPjrUwx2CgMezF7H
8ylzxum7meV+T4JMlT7ptYH1K8nseNq90hfs/MPeJLaLAjERrOy9JP1JlyZ5R5YgF5+4u0lXTQ9Q
qyazT6S1rj4zJPklLI5LNUbQep0mEvsqIai4PD6eTUXWYjCRYO4WPKkJRpZExJp6xW7nS6pWbn3E
HUhpuQ+6dkB55fkOuDBc3UQaXALzOBYcDmu9Fz29fzAB0kfHVRY/fBNHqaRjIZ3W9ncA1sVjJ/Y0
b1ZwFrYGDj4rpPZJ94C0YWjelEDr3oWkX8vmnQA85ivy8ctYE15XBle4l6VzGYy8DGe0JMPQ0KX3
uFAvNn1I0fWTjHeBjPZeov3PsiAFrMX3QA96mtHaZxVTaL8vQpD79ZgKDFC11n2OS6csyPKy5Co6
3/n27+HAm2BwERE0upAFw+cr7kV2sR+whY0kysicj3hTi4ZUwdSzLEMLQclmz2NBEGvOuqGcRtSe
wMEOZylSleLacTekeNeU5SQ77KvHYAgApzhTwnz/E249PDgec9FbRPxqFPqqFN1HjA80+Pa5pQPo
Z0CHG9WfEOMbsNc9jSdRAG0U1zPKMt8rRyZg6YF1TdB/NReIv97ibiElepFCirtlG3f1t5EW1qMH
txJNgK1FZ62/JE3vG/EQPRtNJ7gCfxRB/iRVqXoy7UDy0h3fFoBXzDMbKH8jZDfvxDPndweoB4FI
1JKav5yUGpyOD01TjfgJfSe8AM6t44usZ2s836LFGK2g5ZM/h1szfz4i3C1YT+Ffz1WD7BY178eO
O02+XFFJgFB6+zOU2YUKZKAc40hdXAj/7d2eZPlr5aVw6d7AAJmn2ej0RU8O8xRtQ+shxklikFKd
e7Rx1EGJGE0ekBCNav0g0Vreq7t2uhoIKfnzIVbsHx3KMJ4kPEV4UW3yXTDAW4uHzBuDeivoGrsg
AvfoqJEICfwRAiUVkvF0VSoUYKWBP343Fe14+vsaSN82KkyMMbPRV2/CEFf7ArG9GvuM6SPK8twP
4qemcQSMTir1+v3NuLOs2gLDtyxSU46pytp7k5SEZMlxp+jx7s5c1E742NOpwWbm8EZVpI6567Xf
ZfzS5asVasDkFoyWcqIjfMWY/0KztjRpQKn9nnEDB/GBBuaAYW54NL6vjqO87FqWiypP/xasvsEt
/KVmpUKbxm+3j8hbMLWUs3gNi2wvpO/V4rD2JuQSAWNs/DbpF93TieRKImlSPzLNyDX4yfbN3n6I
4LB4tdQde4P0LhuHacHHa0T+fCISd3QZnuuKPn7yiV7DLpUJTaZdXuDNpRXNnMkfEzrQqcu5rkLo
Z/iaV9iHeUSIhRTp+QLcekDtiMC9Ibl+9EajxlzuMuQh57JYlqwRZL8IpFxreGBAb8j7W6ikuEOD
NkPJoWgpo48mMby+8q7pA51tB3eM0MygOEfFkpSpSAcPjFkVWhrXLHcCLEgjVHyCFVdU/QXpntBK
3S4syjsJdrmdxjMpSRz4byq555w1o9fd1lhsDWEZesoSQ1kknFBIJ23zfOWThUD1hJB1nQ2Gjoep
6bnTtYLnGxLrXLY/1KpWyzVt3nfsSHHDKvZ8Jge5xRazdzw3KnA0HFfAuVQtWYT0xEEg/8xvwu8i
atBpSkwOkuBauC0XaNK9yP7c1O1oblYtwgzB91GU5OZH3ohs+O2xL6b29rSE3iBMYNFlQs2rOFRL
V5OQxkgZyY8RJ4TLEXTvFfO1DB2NDjnQAeZEliQcYSDkdgZ40d1OiDnXqI1J5JHAb2U/kVfeA0ss
MaOCG+J4xCvYMFtubhBcWiYb5xlCd76T3VckU6BlBQ6vH3HTs0azLPNQVyK9XmSUqUEppfe9nfzG
DAFeOlvyT3GiZjQeIzTLSouIt6GVwfBNX2vijhRZRRdcAEx0iHiOS5J+10DC6GI3USDURlg8Rdia
P7HNe7C76tCnJrisbVeWKvBX957PEkQCi6lrEyzzw1KU/SgAIOxSJFo+BrxASLIIxjNOunNC4Dau
K2SC470gkLSPsZVxLcAURmaut7/JiKAF0U/AgtruMmEkTSwvwjRIGTxqKpmderD4tfFOddRP2Egu
G6at7QiuRWHP3tMHZJZEiZtpD0D0tomABwxPM7f57NbzccFXIKDx0KCT1hiYcwEdTpiIypM8ANT5
JjxqtcwUBfHdAyy3hFimv7hh9Xzu3wxqomoQf3zZ3//xqa1VOoONtJcwE+LACiOtsTo+C40iTuz4
jCqQ4PIwnZSryzuVmGZb94EJg2GuWex9mhcANPQQRytyYRWJ4bIE5jqvZ3Gn+X6Q65p9LMSpAFln
m70aMsgffmj86BT/u5osFCs6ARCOvriyM3+g6+V16z8uUa2hBCZPpRnhC3ztgv7PgoZ9NBmluGt1
T395+X1vgzAWaD3SAAM54PIDSKgU+MgPfOcDizKy30z42tDoNydKm9UBYhfhXEiE2Ufk+T9lT0IL
fxHAyBFLRkQITPS/K6R4Wy8KDqVZ75VKGc98hAsKmlBFHvZZrLMnSSPKU7W4orbV9VENRoSRSD5Q
JX4k9Iyt22EVH3hJO3ZnsXS9lmaeQB73x+umS0vHdx+62gLjGXDQETj9H/czIR4U+DQUyubPFfhV
CedjpwHDcewav5q8A8gIyhaR5dldxWUlCIIbqtiSm4y2Hc3C4P0MqVlSeZTjzSKlfXr+100Wss76
xRcaDSNx12JQObFIB5+vdUtgtBVDuoBUDuemgXZvhNdFts2yB5zpQzqZqcQj1R7X+vSwcKByXo7d
Qi6KO9rWz1qvG1qzVTtSyV20efD9QA26SE03LWGhCjeXc35+qgvR2M8KnmbabpW4AbPT5gxmcQUQ
wb6Qm0cNiZOHUH4vgdPOeDgXcz3PWTUq47MZgQ6h61tbv7/Cqs9YwQJZbdW32SqvGwY39FYIiT3t
CijFlG8oRw+kEseqNRkgGjARTmynBRiYM2horgtVzC8SLRfwxyvJYeRKOovkAa87jKrxvPhVUdCV
CHSqBew4UJhzhW0n1F1XPlHWdb0y/cBscG1l5NgtHdg3tu7YLgcREHpPCLKX4zD6Q+G7ehzMWDuF
1IlPtUrGp5lWZVg7Qs7eaWPxylqWvB9yGkMQrs7e5Jlwnww0i4v9qBCwEBHnmzooYhnvzYbid2SK
l4Fd1kVqnupRqsKgmQlLOnwwdjK9KLDqDHW2jVlWvX5H9PQu96x4O7hiAZa6Z2KTKv51BLG6NdCt
4BCndbdYw+oEJGmzePAAgOOuhX80DKHp2BrLMtIVTtsjurOFHrFwVbczt9erWKczLjLDGZRSjxwk
H+7sI5ZzW1Lw+uHrVzh05wccvQ8WN0/ESh2KFJA40QbzJtWfHfqxGjAY6coQ9Kflv+6BOoVQKNWB
M57F5B2KcWzaPJyOzChJHcZPPaa9gjXFPHp7AbKEbXyhc6mFN8y8+09ppkEhcLLlPFEcQV8C+1oK
H9Y6TmvJ0XTTOnNS7Kf5VjBCeNUT88dOWKXmJb8wPRpvvzJa09/XivROrtc78hI11Qc42hDPmkQV
lWcGJ68Du1yiR1OQG51aOagC+BLS54mDvcZRc91ba/dMoJvnBOhQZ54y/XHssCwUwJliS16COycn
01d1qGoCS2M3hMnqvlqlmVdnx6tNoObfAovhQH/E8AEvizoVQxrrmupVsgsJzRP8RzJA1Yj/gu+c
6cvVUpCmPLGiTRijv5vZcc1aSacAHF84TEdk7edoYyXFnHGnqZEYXgcw9StOfBtd2WqAtTL08wan
wg7AYAFqClNXEtRhgguNZMiGKgjo0cWqM74GOhqou1sGNGkW9FFn26lIgy9wqMo0ugLbJdL9OaDN
5/8F9Fi+mozLSnRNVe83Uzdjlv9XEeaEQ+08C4OwtzaUJqvi5KyzDpWOTrvVjITU5AOLr2jjhwRN
38p/hQu2HyB385nTgkmUA+v9f8g/4Df8QDa1ThY0bOpvRI7HbYSJsszK/lqL/oBW7JG3Kprx25nI
VrPlO2GU1hQ2/yBccQD+pwSdytLJhnnyMFDA72QntJcludchvHPeQqoQn1KYDpWFbt+qfrfRtdVM
e+VfDDj1xa0mr8HL7PTdG6vZjqFP/pB/x5NlnCJrfztt2P1QvvwPmhZYD53z+dAgoOL3H0d+KJWj
JKLiCROR/Syexl5kZmjtqQbul2ZS9D0l1DosTML7Jaa6qnFoGQ3eo00Z7aulA3ojoFfKFUpr9Kvj
5pe9DQntREW5FcOw9HnFhLG8y+74nPcwbDfl4jqitX/TOyMacW+qZl3Zs/WszhppsT068nKNIBmN
gFiVKUFOi6s99sKwFPhAHVlHP8b8UB0/VGc0Cl9mfoigMLWoTIeYDycdWdXtBh4VgI47m9aQe5xh
GNa7fDWAs0pFNWMsflqpSSi14oRzQsot0lvgy8fhRxaTQRVwN8rOIbMEkH954tp398rT4ZWaGyak
tINpiLKX3IWRS81+Sp144MPjGv1LQ55Vjc6NskMupqSHaeougoDW0sEBA9oR3+kbbKcvXxM+h/NX
G4Q/TLviF9k0/pR6BZk1IwmO2C6tQv13FguthCpWI5IZEIbLRAbvkd0cS+u1iN1pgyVno5IM2dF4
KckNSdrvhXU8cSXcVx2qKd+3kAwGosdQxHUMzhPOP81j2E0YwExJCTy6ghdVoX883U5RJ6DaeDsE
QRSLW0j2ew2yu42nWCUU6R+VKUkhTn/+ZI9X3yFl21jmwlhXfEqWgfvf8zyvPM3uJufDdCNV69UU
zlwyfUF5FEHRSeWxSg4ctn7hQJdBfKVmACYb6lRktIQXdlwVb+1bdAkyqBVI62U40MJjT4K7RdGa
mups/9X2Rcv4Da44dFVVEzgCjzUaIeJVtisxAT7S2XtKbd7hdGvqvxIYNhv03d1hxDPVjuU+TlPv
Zo28AL0qs2ZKX4lBW8TDF8QhEYQYcX+yDs6IMTsu4YTx88uUtvLUDn1Tihf/FgPOckr8gg3Pvrka
0zdtajsItQ0f9vUlCzQJiCNy3zz4JaQlR+IraVBM/FabZijM3WHbcCp5/j4lvulEUztTn1/KGKGa
QBvcdK2ztRD6BzDfsvMD+YKV2zJBHk7YKajvWvz9aQnUxh7XHBVxN93XWGtPENTCZW+9IZhp61+I
YmXHD7f2U3klgVSFS29D0Q+AbhrPIKMFJ35+BWc6M+9+uDzve4ZpcnWYUZE/D8BPt3FiRA5L7nsv
KteCVWPLdpvfUgmklzDas1AqW8Z9YZJNCPz7HypoLSCVKkZ7tUKueXo9+JQvmi2rYfbmFYBejfjv
vf4FktPch2SC5eU7PchETQ6+lYR+UbI/HyFlRQyBDdqd+d8cEbr1O0j9CSBAM6LwJF5nm0zL6q3Z
F4JioyK4kHKHBkLGud6JsSGQEDrtkTs7KEcbXrsxwPT9Hu1QLvBsLesrJCqjcyz8I3rd9a5DqwiE
5AP5SBv3afzff88P+twWZQbPLWdEKoiH4GG1aqVL8UYnffv4pA0pQMSKEsXOb9FKzp/5KnOF0LRo
Vf4FBDh6hbRYpRVM0my6c0DB+QFj96evNHn9hboIlpj1Bh2TLJV5N7Tlzi7lMbV+dhLKlaR7LXMi
JP8fgEHTLOiQy9CvOwXr3A8tQoJXckdle6Prpw0cJ4qjlIJQFlvmcG7CaeI6kpy342uJ9A6pYKSC
hyXt4DLkO7ioVpz7XUB2Zivi72B0ikAgFbcnxmR7nFNRfIyUqCAbJrOTvFb1w12nGlE+GCNw7TqQ
fzbAcDjC/qYCXOqkMjBdEFNuvDPjwqSYGSSIsd5ryNl7DfCOpDqf1ZJF4gK5Zzo5KZ2wYjVmJCJQ
xW2lAAJFyL1+Mq+bMEIvHeYFL9CJMkowMDiRJvjD8dbOtO0gOTWWLHLFVmzIT8ISOLW1OZ9xv+xJ
n5SiZY0XOZaxAqXtZZGl1XfPLqZax3Z5m+L0683elUEnBC5Pby0sIwx/mYf7FbQPPzcEfV+yx/ae
aTSvKPNq0LYJ8uWrXZq+UEtsSUN+TFZAa7y6DZAGjzKViHohUFHXG50rxbfO/nxN13X+URGu9S/E
KdceBbFhfMRYI5DejZYqzKoZPSaWilrmu5d3mF21eQjBvWJiS4q2rdw9c69mrFK6zmDU723C56sa
TFwqmAxTtvgNEhmvfnI0fTcPVbfFii/TAqbyq2mNoOmxW8Amh/hK5XH0/7jYWDfpUdoyFnbWwGMs
UdQpTveGA7jBKDBorOamOw2uazFF12U6Q5GkCEvVNFgyE9F8XgTU19rLVsnNvxQC8xAEatsCEhqz
s1EdUTiHN9k27Vwvi/GQR26CYN+KPf7+zkIiULU0O8bo/bE1NS7ic7rMaP/9jbOVz0jVntxLoapH
q5u5JvoyQMzkAxsprcmmeS5EMC2HnPQiMeusm4HYF7MSJeokhz5cRr6VbbDDGZJJgGuSHXCiMwgu
x2Eil3WjDNeXuC3Ap/No9qfg3HuIcrV238W1fUPsb2LvGfKddn3ahzariUDIWVU7+YsVlOKkRPxi
tdC7TCs+bXwuKg+ZNDFGTih2lsSVKLCe1f0RUuSOdP99nYoK2XVJet9OmLwYMmR9MulzjmQhA+xL
Rgm5SzzUmDaOKROqaJnu2TUgvX/gdE3HvMQd5ae7W5NgpLhchD5pVN5m4p/wzyjGb6xHj6sajE5o
P3qnT6Y8gyQ0lZnf4XYH/mcHPu2uvQCxkhl6IsV7csWtCQ8MESpTaVgZyrgc++rpLssgnufQhkxj
Dk5AZCzcmDZwlMgWfveiWVoEDlv/OecGOFtsL7clynFkHWzwMqp1RCD4a/wnPilhkEcoDbL5vIp2
4kGcopsOUsX3OXiG22CRF4dbGArS5AaiPHCQX86kZCjIdv4o8mYQkyAsamt6kk0/GqDnXUBDpSPz
Zmd+bFpLMj3ECCELHYd7BLeaH+r0im8326jMuI1svyesYumcExnqKJcDXxsoQ3nOq9vuPC+OJkIW
MnKCFPtMeUXBcY+Rx3pJkdASu1WeCF2qirXL5cgdSJvkm+aV5sA7uc4nJMLBP0EymqBPOF4SCP0Y
zc8EzoSBxgNaElVIBPh2lqRTW+RmOmSVcu2it5xVBX1MbvwGDyBeES7naTf8pVB4gWCZHZaSGR7r
iTcaYnNNvKwdryMPsNXkQ+o31FkdgyL9vZN0/KfBTnvUUaHmBiQXFX/CT1zsBvWAgZ0S2BUSCd9b
nPTT+5GnOPPA/UeGrFM2s9/AVupearHwUFQaPffu9WzBlL6ooXCoAxr71vrTLBJk7taim379DSXO
ptSW1au8ekAmywg1bMim/3Rhy31WAqyKbQN6B+WP99Fwj8RihcSGrd87/oErnnT36JnJJXE+Rkdj
Yaz/B8JZsSrDal94FS3L9Y3+V+VreBG2esugzEgJJvGn+Rh1moXcmhHz+0+ZRSqv3IWanAjb/76v
zjIsnEEPUHgOpOoDPeTSkuiD1oX0RGYxdjJ/t0uBe8HXl5oe3olKwOdvWCshrkJG9dh0chEm9qOt
v4Wcqpd51K7ATmLRBeTJC6hThkDPh8dL1bYHvcE5mbr6BsQcroj98NPH4jvLH4nSC9PWfjXaTlAf
6HxGyB0H1/XpUZD+ANvd62qFVrsp5TsA9gYSwj858dWs+rocSZKRjWpRarwpkfDzU3KhLQNS2r6f
fpK5sB7kp7QjM79vSG0BKsjiu+dIV8qZUGJOzRL8yQxU94s7g+yF0yNIi2FZHHvl+eb/VqqYEhfh
/haepdf20QnBobCQwWbAgBW0FgkPl3Nl6Er7pwU/G2TFZiD0YXp0DH80Jx0h2YyBOFZMw4JGrqN7
G0Jy3YojGviz3tKX/IO8v3F2QOSixRedKC7x1DUvfa6ERB8YO4AweSdvguqfb6I5x/hFFKWQna4i
aIB1jk8SNl0cTsWdyopBBzOCkh3Fm/D9ixvbT3j0pWklqBIM0ATmQgU4QQ62AxJriltjTfozQm+h
OCPplq8i9YP39xAMwGTqBciQYX6+x71lE9hOKNLWlv9y+bRvIgKWkGckRjs5JopitTrQxR8X+fcB
ameC0JN2pflhmIUZDcdlWZX58bKLbOAgDYzn+yJ4E93WZtUaLJk2FymG8Bn/OvAwWzb37s9ig2ph
fvfYN4P+NvhD+hZIqEvVZOd+Hu8P/ALN2VJ+5mrsuoajpS6pzIiXxIVS9XZpkli9UkULw6x6A7zE
flHnM+y2TYXgpkIhkR22GeEzJePhTwtN/H5Dne/CSfOFCEnoccGpyyIzub8HyBdNObBcHWZ8lhWz
kiyTGp2qOD/SxWSTcXmYhXLkQfiih+niLSvU2zAg62JZxSTbMFwUfMJ0DuNfHCC+KgFH/sqstu7C
BS7T35EeELsH7Sz9q4ix7JXkVk0H510XWGerzJJgB3uShErie26ULCMGIWOSE/91peGK8eNYgvDN
XWpoErkaOfaKEx0f8XUE45q5upPhq39yWQ/K2FHwka5DMXCwPC5j9TDjjGm0RzHNOfulerzkvbs5
Ex5+RxSkXitFdqJTkNTdWq2tMEroXuofhZafgBkXiFKgvlBChF+J32qp3brHlJtmsR1nmj8lS9wP
UtxlNkRkEgZ2Gv763rK1MhCPej8CLRsKa2zM/TyKCaU5Y+QKn+bg1DpwPTtccgLRneUI3fReB4I7
bAuXVfNzppZRUOBD+N7L9aGOlNzZjY4+H4I9W7A8iCOwYmLxn47fRSyAVmlKfVJPIhdC00ofxpYH
kciyJzPiFWrLyLH/rEOQmXjTUuNrlnnOFy0JGqFtG/rRH6VsMx7u/ZAC7dBQl9j3D5I7Jjl5Epxb
tFiPPPobku7r4IxwSTkYR7xfhF/FHe/sDTrwTA3mDzQ3l2WtOAiLPNAsv5xS4Mp2RhlR1lsVRcbB
1m2Hf13owfLW5A2CTUoQDxTjdy4+X9rTsjZhAp6r5xwZYVkS0kTXGN2bw8Sj5+93m9rOpSZhsPc1
LbkjihsB62r3EyXUxFp6c0nHUPwdSWAsd5ZgIKW1bxrxmEvVjO3SUFH1lek+bbt6WlNzyTu8DKzM
D2Mbnx5Un861nvvFZITeeWTiF1+kFnGvmAuAm9th3tnu2BjN1rT+RAz8t9W59ajEcH7r1BECLdM8
MnArh6cXyasl+K2c06HCJbSU5ZkP/4XpRABtbIqx7JQVAcXyvAre6CNimMBDfiSPhA/Q8WN+84XT
Csv0Iv22PtwWnhc8VDe0yryzbjILx6FPFzQ4qzeLioqZbpYz1eIfRoyFBrDxzmSzx0f1OpPtmJ35
F63UFfiAExPlF30GtaSt8lxw+6uvfuQk1JhTXjR3K4ij77U82NjWa2fjZwiuUDKVHcHeQVDG+KPH
WBb/Zl+2OMOZBYV0BfiUo1asBjdaq1F2oq/v9OLJ78uQn/CFNbZ/1iK4l5A5SkNDjPNm0xlt34Ir
MMi0xr6cMUgwMlKtlGExjywQBuTqtU+wAcv5/Q+rVQI1+XOuSNqm0T98/EC/cqQqROyK44rDfEVW
w7sU1DPmTnM5TYs7kIPMP9BTSa9d6TIGIs0ydRKuTPlswApk3AM1vl1g9dvD835tfQXtv417e3cQ
Barj3rx+eew0fg9FCXIYPUY+5TKykBaIgxVEJJ4s0SEQUg3GsyD7XuIhwlpVJT7b/s+oRW5QgxAP
36slkIxXy+8xZO7+JssxRvRW6HlBd7GFfWad1VpTdwp6vo/5IlP0HuzCljZ6kfdc6hdbVgRcDqbW
/MdcZDE7Et6Nt3VWBhckXRCPRu4H4HIQxzVEK27p53c2il4QJCFikkL1p8WR1Bm4pmpUh0xNF3zg
5Ig3ArH8iqcZgSGmdqdFGpl05PaJarbus4RGDili142Ap41qJ8Euayi7MVkX6MIVCAbLioWYdo+h
vgk4fnnCWdXYOJIOFYB263jGwNgAQXz54B6wSU2wcEr5INab4vX7MDDtCXqs3rPnQy4sU9g+Tq2K
pz0g/V3Rqfcd4tuC9KY8sJ/vr9fWvQ/eXZjSl9z7hayhVqommaPRyfR9+hD0FHegEfY8xrOjO/zY
2OPSFDEvwfa8zHni7X8EWmYcrIL2ROTvGX8AaG3j+L71SRD6LItFC6AmZZik6XnBs+sMoLoV0xyS
UZ0GTf/geIa9grFXatdEai0byBj7fsemtm3zjWCErXrW3X8ohc3wY6WecPnqrMaLFPRgcK5BIMaf
Cw7Tb67tDyJ5up6XxV1HA0Rw4TpfL9GlmB8Axlo4/m2Zu4nwT8ghoqj8UcGmTGc8QJEPs4tC40iX
hIA5jbPy7rfaECXledyQeLQ3IgsnI8u0DWt/I5Yd2ZZB+X0aCgFxy/SzlGewxWsAP80hl92l0K3E
io1u1Oq3r9ygZzanYsfHX9T3Ps0iEviLuXHTvx+AALPy53SZ0BPc4ZTRxFrM/fnGjui8dZo9ybgO
V5EOohEzSspGo2DuhySSKz+SttMALF94kUHN08k+UAJ//tJHJrsB+itaWDkopNQkID+aKIg/uCQI
idw7LPqN0RUh2NZ1JHymJLRt8eXGg3nTf6nRHrJ4L13DPjZkgpzsfe8Srj2iWSPQOzEt7sySLaJQ
BVw5vzBWpaNx7yoel9X0s7LlqAmGObVy6/VGmY8bNbkf3HAHbOAci8cdmLxDarK9p6EUnX2VyNDF
UjoacUInVEXGRPuG/7ywJSGVL+SA4hAwt9b7SivdSPhTYZCN3GffFANDP74oNmCJYMFSeJ84W1FI
0f9OD4s5qn7zy7CW+ehU2uAqlViwe/SC4+tfHzBSg91PR/RNzGa2LwQRf7QHJJ7u7uFQM0s/k/3m
v3vzHGD+ebEdlQS+h+OgHJR+jFUE0g1Fx85GpXXlNeOJO+AnHfAOZ4K5v7aXcYmSH+Oc8MU+m+61
GBMtXtXrzY25uCW2344tsaPgT/TqoEOgfHnY+/1jPkSmiLvk2Wm54tt2Lq1PS46Lf7UVNk2G4kaX
hogATZsJwOnNyT1XglkkbcG5Ixp2XYe9xOv70IY42zvwsdw4qz3V0oroZH/7T2l3S1fDBsQiX2CJ
qdO9r/7ehrrdLRjLotVH1Nh//3EzloaBMCqO0xY4Mih9Ol3CXtqaULiwNdx81BwYriT+Umj0X0FJ
wcSgMOJQjcgbKY3RFBdJOVgUQ0PvTXCY/UI2ydd+bwAS9YtKdR5zxMYDlQIhYUVIUqKJCX6qABDs
qz8zsMVuy53M2mA+ygquUJU6YewKHKRyulZ5ZIlAfh+mCYajOFtmZSKM+jh3RQCHmOC6QrcL0Edu
bLt40ROrt0QkEIyLjIuAYxMxsMIb0fNy5tIhkEiP4VFPpMJaKvJ+N4a4TBBlw/NG8Nx5ShzwEgVG
SwGpX/vOaYSFVoyh+9XgMgz5C9lFnWIY8cTaCY1MqYwkzlJptU7pJ82uyABpXMmDAvvHEsrgbTeo
5boJigIr41d66iZbs1oe1eKc/JKBICGDV1SiB+Ctu0NJ5XYV4bdSshM4Ro63HMfk1+VBOB95rsni
THmZeU72e62m2ny5UsqrxumIQgMJvbVMm1XB43T0zw3t9ftP/sZYvHVrx8zenyEwQxgsRvyoc+fS
kfZG1IUi88XJKtW5EUkjFF+uUPtka2mCQrmHfdZ9aIOO/OeOMQC7yB6zpKE1wdfMgdB5HqP73wzS
F3t+fAPssaVfn8cqSLpQNIBdsob2EoW3vAx6q1yv/HUjPqUfdxh98X+w+1hp5Sv5WgFrYYf3OWTC
NCaDcY2Y5GehRpKaPNDNN1Wn7KzcKLe3jbWg5RPZXLnCNxeeXi/ewd+ORnH8aBrvh5aCipAjhB66
bpZB3z9MxLAm0T3srx0edOif3pwoEd+5k3BkFAynVmUqRC1DkL+GTe7eo3HDslTS6a84Lg5TsXlW
7gY7W3u/Xgy8UbuGhDs8bt4PRRmUfs0ZBswE1Y1lRAg1cRcRlfimwAFZMZXJ9JAmQUlLk2T6Vm58
py1jcytVxULPvOuRs2NS04svz1sku80+QwqWesy9VJbHh786JGJmcWMynzMb8eBCuwRtHtLOWwI3
fDaktzUzp9zGo3Bl0rkXhWRqDjpmlKxKfq8DirQjX9XjYmBdbkuzwijJNAsKaZww4GYx1PLkNmc8
Ww1YYi+rVnQVf6OJEPewWjpeNpCjSmHA2BqIesRZDM5bbaUz/mgwW3rv9AbQouCIZZzlZi+tyN3u
j/atkrGEUKf7r9Z7+hHbeHPBreztzpH4NwFvF7HSvucL0u+HaxQgm0JGJHsOUv6Z2dOOBP5ngrxf
DMlCnkEx75w+IBd1JJ7lkz7a8TQtSoqnSvrbrKcR84s3x0MeSOA1jwxvCbaw58bVmqcBTqWJvYn+
iVT9O8GNfa7xvVtexPMEKItR8eE2DvHephHcGToYuP1D4yTSv3oWkQ762QRUUbkBtSl+7g5E5bKG
/UwKV8K4f7mf5XOcvRUaqYyQN6z++33i7pNb1yUrICjGxkFBu2r6L+ClVCsatax3q1qf4f6A8f71
EwYEl7b71/nTSndfFLnOnYHltFAOd+DN0Uij7NVLB9f40lKVsrGbqRb8ql+TGsq/fM/AiiZR6fNP
V+8pnLCLMBKKlPHZFOhpkiKeDWy9ndYuazy+2ptUe6pjBEys//TICxOglLIQ2L+Pz1273ozNybXV
jQKjAfjd0iY19SYi2heTzf0RZKJsZbo6sZI+CKble2X5ICZYlqS0nd7n43m31S8sxJ+2dF7hNARE
uyhvEwAKBAFxGJmKpEIi5ucpXpxTYiQUquUqELkC77DKnD2fu36Av/YdOJyh0oy8wCx+Km7Cf2xt
gqm1pMdNTgnq3P1IsM5A4OFpZeVKMU9M3Z46gPUnDGq/A6odK/QsFX0msNj6PP8zWUzcQ+bRjR4k
jbv7VGNzLRCzl3ZDLYJi6r0FpwpXF5i8kcItfj5B5edhCNFvdl4DF4p96jf4Q3Jw78FrirJjd+fe
DpMqbBKaezFMWNYwnt0z7CwKpKALlVYs8B3ZIdCGxXF6J/zPtLGpe9e5QElLs7aeZsVOx3W1am6j
PXUd8I5izsUoP9lOe3RZEQWzOlAPB5plny56PXWzrqpkvX6nzbBz5l6M0GqxfpayVJNDJSM/zU3L
pO1PbhapEXra4w4z1GLKCvwSA0Ync951nLFsMWVk8ehiW58Gie2ZumN77Nx4pqakdczWwStC7czh
0H+Nj/bQQIsXZw6kvj1r36igKAsWAfjNU5FTWXOX5WZnyIHLRGTmwiYbPuR+oM8MdgOu6WqcRXkK
K5eauHFk3tyYzzV8Zg7ubVJJUGV8iDRLGk+v0K/beC8oVt/BCLyteXsW8Gj8PeqHkT4DN2OKm+YI
VfEoeLpliJDvtX3EY86xUIYXCPPk3+LeidAqrbDGO7YB/Lq069o3FRSn2OPK4SIRi060z0iq/kYa
TRGizA7eJqkI4fpdbDCMwAE00YQa1dFGmBKzyUxTLGwvQmU9zHUiV2sod2JhBzl5MTp5phWryldZ
zgxQU+pNZYT8R8D3YczN18a+592i/Rcs77Dwo6myiHoP3t/FlI9D1q8LyO+QyYILHLLjgMXW75O1
rX0UzVcv3+3jT3AMSBAmkbn2zKmP7mp55l3sZhXuvZ5Y8aUUjP+DjPiWgjfcySGN1eRKoa0zckMt
dVMkUmThLWM9gli+R6z6633Gj5TIsjgwl5iZsYFVOHnSi5uo1wbNR8OSpTQXtFXiwIPCP80oX0tZ
2aEYix/nETrbYcZ5vxGcY29QvaPa7B9Q0RAiiEHnFunEB1JAas8I3fOPvmiGWkoEe8IcG0TysQJo
72MSFw3DhCJT0l6N7KWdRIJ3AAEOrGiVsIehhKBwFU6Ay+X3Jv8r/akesTZjPVCy0RWboJRjNehU
HjIAwp6KFXV6fz6DFUcIDBff1vSeox6sBpP13AyJMaJ/u4acHX+mVp5qQ75kmjy1rN2VaoHf05/b
2OFRaknszLESr4J7ucPCxVoH21dQY4OXFs5x0vneNn9xBhBn6eC1jO2RYVGsBmwaa1wYaeqTaHzh
x6yXF5V5e75l9Np9SlYge8kHstEGCgVZnsyMn9hlh99pX8ZpBJ54GgiAtUEQJ6aj+EfjPrgJwUCt
1gQDaLWlSU6lZR9yDj24ArdiTN96xJQdh2R2hZknNeZfCNn/jW+NHbk85OWUjFFZXZxZkAfirEGB
TkhCbVfWqi2vrGbTphk4xY9N47x9EEDz0Mc4QT0EoszWJOtzwNxud/tz13ETUn2ZHUOPphKQJp8p
dc46gLY9PFXtV2Egp6lJME8Urxm10W8N3XW1itjdYu5it3oJDXYdbgVoWxMm+uJdV7WDF8Nl6wiT
RyIvVj9UAfw4zm9vFvDgafgviwYmgr6b655y3N9wcDGLku39RfHoacU5tSWbQ0jBbaFpmGh6WWcO
95Y8y/7XHGFpi6Xmfh22pz5HHvgu4m6dR1sWI4QenwZb/2c7C9GUS9v1m70cQmWrlQTR9ULWo2Zk
WcPWv+l1T+QEyMkSpGlLLV6lWx3jKMccny7rGDIEApct8cQLNJBgzCFX2Tg8YyBhWa2ok/QYAKlK
/1ayDMit+otksqs0FtbERhFJuTVGo/QFNpm64G5uAEx/0IJhFmZN9s85R85lX+cnsI+4w5O8RODC
5RB/9Ks9JL0i+PXypu+kqbTS+gcmyI9ugX3VqcRzNZbp9kFFeUGNFrNAtbJRojwuhRtmFTNWJsuW
bFDLSavMXRC0/HEEI+xCtqVyucI1E8F/hlY9uUGAO7LdMr0NtapnYkMFDSss6jHsbxcYcOquKpWD
VOJ9Fx0rT41mAG8CGeVKdtIEwJi/2WNJASiI/7dy+5lfkYkOg3ED9InFZRl7Sjg+8JHpu+TB/leS
Kx/OKn5C9001qEsxaQatcUk4/Q46qKjeL+BG7wNh7IpDchAOxv1DB92Qcr//nk4F0FjqRM9rD8wi
M9VTy/6L/QStFXbX96y6Dv0qLZuUuA1uLSGi7DKZOBFz92kZ1xvyhMP7bRwvIpX6i+5qWCIax7Zj
VgA3A501Nn9o91Q56wBIXrnDsgPWKxMx1ZkWm9XLMXu+hOiZdvqLJumntuyG0A/hrTGOTPnY8W5P
6cjyUKOIIZsYTQboRxGzQhXqKfTxAKvNOsFOEZkypYT1ZtJpcAJuZM249Gnc+1Kx4dbx6+P1yHUt
75lRdTP2P8sc8aqnWuUSYQhUHehjLBGiPj+QAv/V2bNBibngZQEG4+mkNTe2LDodmf+IpWmkmuWL
+VDs6KIp8/+0WXxIcr89bA67wAmQmj0er5Jrrwez/UsuRlTa/UJdfPRtdvM+qjilw14Hj5FePvAl
plOzmDeP+c+blk6u2UzIg/Slgsy3b/Q7aTyeNikYpIR9CrOOHLzxJCTz8u0DXZQpQHNkKSYaXQa8
5DMxCbgYCf1PnlwonWKeckdC0khgzHSU0OaqaS7Hza2FzN8mug14GCx/2qa5UClz72AEH3EzUv9m
FnaZ3QYhE1yt40SLhOh/vXVwpXMANbmh2YGnhZbBF7PtRZjP9aqlUWjKPsT7Yajr5oZU3ZuYShoA
qudt2T/QTFMbBOddbp0O8wgMNDxnDcnsBULC712qyLY02A5Z10spH3dXV++mLCHm1H8JEA6/3Itn
Ot5dkk3Cum90SHYgT4600x9WQaknb6AdjMKdQi1ptpjuWtmXvMFyEuZXYv0MoP2t6KPLAyEfZDdl
/T/jISXXdMSkRT/FBajU8aP91GJ3OrlLmHRhPqVhsPzGq32b44EO6VeWt3pUraOpVEHRw6ydgKpd
P5Ytj3WPL9cMY87LAmMnPebP9FUjw6qnVcHlloKhzWii0HR2FP2fhVZu+k/4VEamKs4Ek/n6F66/
LlricAr5XQ9ry7I5R29pNWHqr0WCaK9yDBUtY1GOGakbaVUk2YdylDtZW1Is5XnPsLzue1+DU7Cg
0WynF1llSTyKfl+eHIMiZqSWLa3wtXLRAXOuEQUSI29lxJorGvXTILCadr+H2eYA8EavQ6B8KpXn
ahWzruAYSLPr2WY0LGuSEKWJwL8pLmPLhHs7uQgDwXAXE0vg2F0W8PphRoZz6eEHqElDlnwTO4MT
d2nA4wgcSATjOyBjWoNfELI9T7qZTZ/LPqJBPtsWjkJeOQ99RM3zOCO0+dbhdAZGS6J3C2hc+5wG
Y5KlhYKWuPB3uH7+Ie5jr22dXizbVPZ8c026TdciwwjuJOpEibyHP3XJ27aQTy27Ym4vYRHlXKwD
7QarGcBKkUe6uSohERpTcGrTrBwO+JlBadnkGs73nGRHG2ayyRonL0gEyVashjCurd0V/mBuRZZs
E/+1jbl3ZDfw9eGvKh5s5N2QB80Dqn3fSNBBn0HIBr2aCWav7fE+QcQdJlYrE5wm0HQedcpz3Rsl
F2+42CCyScVygWYySIEg0TyUPmls15fFkW2XTFDewgUvJq1mQkWXsyPZWhnLNTVBfRLBgjdCbrjA
EI1sAIIWIMDTbMCGD/rrOq0UfR0lzOcNb4Z+tkE1VhPbm8lU9d7wOk0GQKUSqH81r5nFuuAa2Mrr
5B4Ttanapm0Ra3daZwMpcTYQeKUXUYRvcSHruA4C6qMy0tiB9AT1COYAIRnNs68T5vKVstQ2TYxk
JetzReW8OxB7DivcF+RGWUCaecuYzKfk3PCCtb0EYrZi257Sz6D3x1N46QeQ4NGWqRirVCLmN33k
m/aMdGBkCqyX0aB6EEFzWbiXQXbHW0Ja8mNDjfNP2EGr0FchqDAIgO81E2hSNM21aLNot6UOyST1
EZnIdwXXy070RG4imEVHyyP2PZCQ/ckyAoLiHRoIvfwLoR11ywZBQMT01NsTzc5T3GdrzVXp7Vh7
RwGM7zpL/Z+TEVDfx7CNXfIQwWqZBaIG1xwr1ydAJU2xIUxiiNXZ4IJeZVQz00vh4BfBozUc5LmV
kk1+LGkGgbEZdf4+WN4NaM0wBBr/kPML4Gk+ZmzoIm72DyRHpicCTSa/BPJ4U+0kLRgJwy+gFiR/
z4lzKtEZzsjTDHkHXgoAjKtMutN/W64QKOmnxG4z2TomkCjCy+M8JIIeEc4yFXlYyqSugNDIwWYk
iglQ6s3+8hz0Bv6RvPW5G243VxXH6htc1RbKDipbVeGpI3sf0PdKZuBQD6+z2UWYktbPRM2sVYy1
SN9KqJ1zXQuitokyfogUnRaH0NTrhxZe3dc+JvAQ6p4uwvRF5pIjsI3ewB7CHgUN3HBeJvGOXrsC
crjj3IXMNkpccsjBh1XiEOEoSaV3nF/8XHMmMsNFetQkYvBvRLeZS6Gx6QmdL9geFIm6pdzVqyG/
LDIeb4PwA+FMeHODi5mAZD9Hdc7ebRI6Uu6wnL+YgeivTz2UFynz4shOemDscwDozFKwxmWKdcVj
0WakpGs7wb/KxbYL6aNHA1fGKLf59xvgFkzhPeReurs3zGy5WGrE5cGV7Hd+MtpaT/remTwCk8aQ
RjvPy/f8El1o2df2m7/jR7AIAzfObCIKQL8r0nds/XOivSjl5Lt6uGdRc1cR/SyHRN8sO2uHakgu
CmAAeaBJwNHeIzxgVJ/ehnk2z+QEuddnr062C6ZOE5AUq9IWXnJB9YkQCxDx3ZVW52cwj7oEUSxI
UYZpoVql0BdsBZ0plx9ey+Hx8vHEzVrAkJi6StLusq8YihnIezithXO0+xaxmSY8jJtL1gfjRWgU
myORl1K1XRK3XYhcuwby18cX2+adIFEHX+8CuaqDwKXqijckuZjbtrmTnmxOKjKCZmTX8QtuyOSL
KyOW/+xrDVJALPRo/Vb5/QH0GU37avRqO7aZath1jKsDi/1QYeCVd2JiIiY5jAKhlNUg8Jc0+LBK
rH6FQPtB3YTvPRCt5/PKFJCb/OIId7IWnaL5OYQ6fE2CdaSAUsVu50RPQ2atvTZpzm9EXBDg+AG5
kiErMQJrHk1Vr4jZz5rmhDT3tHvKXX3W7GiNKnuCnEVKEAAsqmMeJF4obVabX7yGaB1EzXJJyTrq
PugFDkIcxHUjv4uLg4b/R1bHaIw0rUKFCGC1i4cYLsAKRbx745/Neh0rVxHKPMOP2+pPzRWw5KSI
o1Mz+85KxRBxs8zfBEB4GPxyKW1QxB5IVQ4V8OK85Fp1Vg3sVkKsI0srVU4Adp/ArpIOo5Yed/pW
0kAsQ/UZn8+Dvv64klUNzlkXlWZjj6j1o7X/dUlBIwxqRwy+kyhUIMT+vLNJBhIvuMpZG4EwGkdo
DMmuc4sxAIlwvFnlTETdUi10+Q1UQBgyDWwXrQH4+trf4YaAttrBMdrK3uUWMtEiF7i1wPkcHkOn
WByMtcksly0mkFc4K0Du0+wHAHz6+5TpLNL9WE9pSAIZ/jA3RACLgyKoiVsrGl/xxwjrueB2P3KB
iPNtBHNID65JN+DMydzhQRDh8KOOg5FCm8tBjLNQs/l3cVxEKYI4xiIVoI1tjboDL16KJIJrE/Yj
WCw1VJrGrfnp0xzFUdhMi/xp+HLjS3sz1pd6IkzgQr4OpO2aqCDAz68QyGx6MDnP93It2M7UsbF3
XZw0RghgNX8vV5bNItorGuF/A3OG+Zi/LF6UW21CK9lTTJ9z9bmQalxUc7fJcxT4fqDhPFi6VkyV
4lVtYNLFrzIX7yX2A58hWTc5W9a0GUCd8ywwVebcfuXUyPm9KtbgiQd0H0M95lBB5WLiu4cySy6W
hqKWY9M3rEfXkgKYcN8/6N7KS8HNxFAgehHgIN6iVe9sE1NZqWMiQQWt5qPFS6+JPY5WSuOfbENx
/zaKxn4/GQQuhlTC7rFgITr6X/no9Pr6ulrz6r1w/NLIOjazngqe8t6oyZiXCj1Jy7tCvP11+JGJ
5q+FZQkoOK0pUQSfAJ6TQ4KNGB6YofwaA0DjhKVricXEKd8NsSHnU34OQcKPAIrZxCY+0qhiopCK
uuiVYkrOnRulyTS8YnWLbOt3c1hTkIjttCGItRXShuf0SvjxrEUwZVyXX+LUlmeEI6PhKAQCs4jg
PBs+FXAU7/B8ZqlqRHSYySA8dMcNVBZEqXP5Lhz7NpowkK9vtYJXI1VlEoCZMoMkNz8XrI1+mfmn
JqRUZlMG4QQW1YK1XIc3N8gchT/kij6kK5dyGLInZwFglLrl0sowgICx/wkydl113HzXnYA4tHBh
g14N0ExyfN9c96zTK8THMo8YOzCrEEG6ZTmT+CGUv8t8bp9PEcRLym1c4mgyD8ipHmqu4yDeEdSD
dxqVvCi8fY1qv/hhYaqmzfymuzkOs2rmU5WyyrrwyBI2bwPcuBnX+/awdQaLQsFpklWyRZLFTt4X
EewDW0GrqM3GldZzr4ptjafp0UNDLdtEosWYh1x9h2amJIadLkw3DuCyqc5geAyPfIFHgeNXGadx
SG6x6ZZQjw5MnikuF2mGvPkw4DST+i6ma1/mIW6e5j6jYqBkA2ih0Olxb1B5T7MFXYtBZstcUBr0
YfPmxGqudWK5BhwJxQW0ARQAVHkMvN8adwlzAFLrcQ+evLOFFiUFC6GASgzkSOUAeb0ig3/0vTWq
jToYkkbQlaCoWk1PyRXZsbJgfdv+tQEA4ZYeb2bo4BlCSY0VzU07ugZ31H4iWjEkYogFH3AgJ1CP
Az6K1VfOSpapyjXtpQY/FWbd2rU4e+U6vEsHAW6A8rawxC1prT4xhLbMH9QAhfV2SsiJGtdv5yOh
Xr9FZ15RRmCqLwwsWHGQAoMBbSX6pIHcyVK/ucDTmbLRWA50R0O5puKhzqNzx4qEx6MfOFOr+qln
RkAqf/+xhWJK8TauI5E68eQqZeqIVT/hfMQyP7dOyJJZ3VbOS2Kmv7FkagpVjsOLphqrJopvpNwg
ao1Mcha+QiL+V6+TFzz39y7ES3rogOfMQ/6vzkSTU2HJfJMa9d76yJhwKXAF2tTJ71p1U7Yx5JO8
9srYDnK1I4zGEDIiwKbQ8kGirQNvbUx8iRrhKIaFX0SVZReee+KdTU3cHqQA02AXPLxGWiWM7Rcy
2DmWTkGSFSHwYzC3U1+Mxl0d/7DZs581ax0wp/na/LoMRAjUMdwYBF4d4Zb2o5DtLG179hi05h3N
LSKLhNg4s0Nq7L822wxRKuNHNHZgccRGVh3yKKJvnSPqWoOqFMnc+b3Z7yUYYk77kj9JjWPiZIPc
fkJNVsS6M1Hhj26KTQPKQ4jkq4KcQeYqscBw2HZ3F5jmlndIoWcbCvAYxefGuHE/1rD4FlSYfWAA
vQ17CDOjKm7BYvVFQXImbmRQs2tCDkR3WtmpWb9nlP9cf4tTT1HTDCgee/KxIQkugINAM7j+N2gK
i47Fr7MRx3LnsqvoIfUI7Fxd8NfqfrF0EzXH0XHtW8cqPe0bNh81fspLG3POoDJXd5dwNUCakoux
SCK2nOBNP/7F+OcDN5tK073vSs5Wb0TgyhyuTioNFfkjYxMrsOS10V23tDiQzo6OEGUbpiJoG03q
XJMgU4eUfQj8HulJDaoAKRqy3RRxKOSk0NRVcKpzjNJS0EC2FSWvn30AZJACc72dH+3+d9pAidHC
Td6n+akt/IdPogVqwTi0mjgOGx9TJ0rV/T6kS3bpX/OHKVRqYEwipf0QuPgXdAycmZfwBCz4xoQo
gXUY3JZml9F/ygm54wRmwb/1fAdv3uuBOXZYGEVma7vhjb1eXBLwvqXFk3WlTd+V7ctZxjtDG/qK
zlsIDHfLY7WFVmsu9kLUDfZ85Zc52Ot9u9xNt/da5yYbEKSGhhUDLa51rM0xscdkM7QuhrVlGL9e
F9aQzCANjCQFcKb/hQMEmnY23ozFI5DZApAqpw26k07WtP3IoqwZZEFvQog6bC0hISHlUlM3wmYT
iRNaGs3M2molVFsf29t8BNyLTRc05MtEk4TL/5QvUBPawOUDFxtdsSeGZnHGcR/uTOrk2djuJSYi
XvSl7IECsUi7Mm5+oRN1Qwet+2kKgKVxt1lYPhoc5sXtJI8QxDGf9XyqD3U75+ejV1e/Ze26Md1V
KClREceM+7g7Q8c5lmxkrv3bfzBVXn+zfJelWZtfWGAFcF0YX5bUOWWgbjL2WDneMzt044PoVfsz
5hFOoGGMtaCwGV2f6MPUtw0S8zOXj6P+24iDRthK6WeAvlcnfB62A3FoomQumthIp7OeiH5jl2es
Yed38SviPkuznzPJq7bi8Nd62UR13CENF/mVUWlv5MvmFJnU6pbKWvfxGhAcNNaxASfDYerhCHUB
sag8V/YbrWTGYRKV7ddBcIKhWij6pQCegjbqjxswOMuqEOaJlrBqZm7fnCYcOgUT6kxcIxYBwsWc
4JuNSx3GtFwOeSUe1YtbOYLhwQ5JiiGoVEWclzgDQiSElSuiEL1PQrz+upIJMEnN1jeuiWVkUcLS
Pao70Ny8tsErHAF0r0lzLknAj+A7R+A6+1X/oJkayAyXl0BlCixawZIDTSHtKtnst6KJ2TzcK+qw
B2E/DFHCaHumV4HWJr+mkEK6QhK5+xviuzeY4f2zO+XjBOtzYMWub7N0fzTApZ5l9M9Df6G+LLVA
AE5tvX1NSRqJRS7F8cFWx4wLJKCb+aDBtie0nFnnv7JCs0aGbpWzWUCfF4TYl8l7Y/51HeaYB3eA
mucpxNwEVJYJUXJzADY9rjU6qluzhQpL0Pm9qNFUs/KJGmEdj0+y2etobKV1i8V1i5aWWqjPLM6H
BWvjq1FRlvmBvbezJQn5UiIltfSz0K4eflaD/Yfff73TMHfnkCNybq9U7HzIhYhS5fCQU7hD2vlB
HtXQCCwiS1TbeOwnMX8/z2epZ6gTuHbNpfYKmabc+SXc6m/MI8dcw+DGykBdOnvjlDrcM07+DheB
IP+LPdy3XftfXt2XDZalvdqSpF4AO1LbnF7oDxpZwLjtlsQtf24xUDpLnGXso6w4B2vrGj9n0Qwg
YqONZVfYJody0ZNB1yLGPX5n5mUwnCkbBUsntO/EcLaoBsT2QQM2zjZdiE/OU277AZbSPQE4xfch
DyeojR5EraV15QqkEJwDgGQbwTdNPNZly1N69erb2lyh0/U+ZuULzsZL2ViDJU6CdIYBMZaMNPAi
eFtZpaw+/2ugt7wprdhEMStBkLH0q1sMEqVFOcwI0gzS0E8vRmyeha0y/5DWQx+BJFPD9kUVOefg
Ph8Zf05zZcAb9XP8aGpopBA79nO1vmQ3RwJkx+2T1GVUPOJf3WKC0uIBdff/hhckkqvKTeU3jHXK
tIoNw35EVC+RChQnpG7AycrIHGZWSyqyS34Ynhwt/QG1k4zM9ZSWDcpwA4lGXffFYTMb/shA/4Rn
QllXRadSeSMPC+ZlOn/t0r3uv3N5nOS7ss6aWAtRLPlTeOoCcEdR06Ee5zj6yscNJssDFkGQhy6l
GVcS6XqtTKWOWi6vfBkj8jhqkuf+cmWwzJ/Ed28cNW0OMlUhr8lHNLOTdSG2W7qMwG2k/D/9QOJb
SszU9h+qUCRt0hPKyqNAGwdMJwpP2EFX+5rXhaPemOXOMeGpOv+Y6FDoL1KIyppRP874Y46Q6tm4
FRMqrHWEDt91Kz2LN39/B06LrHM8lI5ybPGUiEWERpI8MmVXIvMrhrEpdPT3S3AFNWI02RicDgUf
x8yaQPMXT9o4Fx3FyNB+TI0E7wqLcmp6ZsCbVK2opvFeC5w8scU0qLGaErjlRBQE4+gwu8oT1apG
2UVemtJHTWmtzT2uOcCfI0EcbWij16JNZF2pCQKiwFqpmspAN8OELJgoucTzIEGgXG76NSZhB4ew
jrbF+PwctJx1jB5KwywQPbFR3cc1TEKFrjg1eTKxN8XLvnMSEEwuxKwraO2vW0px5eizs+WUqbeX
ZZoUjpgkZYCtxbfRx5RzLT1hQKAzSzBknShqIsuELUaDOiZkt93H+9FkQ//CwEG8nVDxjtGkJTFG
IAGgK/OQwZbjJduJBc4W89jtTXGCztzeMfMLyXP9pK/knEOAsf/OWO56LvdtTy1VsyE++7RMZckh
oCf6qoXI+7diOWLYQpLfMxtbUCPnkpBVFi68Sbg0Wh0dG/eVP0O02p3B6muucuLZD7n44VmrC7P+
W/jzcRsTgy+FHLMmGK4Cp2QHSLbIaZr6iRrt1RgK3uAu40QgieK4+gebO/7ifHx8huofFaFxbPAA
YB0kHAp9jdzwC5+Lz8UFo9UVp0dExiDYDa8K25gfPMUqkjfOUiopz/ZJiBj8SKvON86mXGA8lX2+
V6QTHhr5VLwNClyTkmfqHCCJzdqyW+Nkou3tyY8voF1q6Br8DsJm/s71gbNRRRBwUb87K8ASZV2z
5l4v8iWf3mfXlvPJyH4czOrkt+3l8rAWWtB8wFk9ROQDBjkKgH++IZy6Cq3bLz2X5fKVhpXK2Quo
Lz5opGxbd9I4nPLR4KONuUKLhkS/aD6yQj8gzjUSmYuOC3LJGzdj5OwYfPCIyYwUU2u1tpJTJpRt
YfXfV11T2k5TQq6Yc0MA2T3s3kkUbNEKOZdoFzErGp4PvVXEH7XAclDVytVOeDRrwN4MvJUZiWtt
Yb+/DHL0tMxyo+CelNJZlQQ3v3pvtcMTfzTPoTks6X59e1i4fIXtpnCdgW4fihgkN3gKTPkax5of
xw/ftyydlIY3MmrO9Ub2ExP1sGwSeuTNcv85LErBprKzJVGzrJdkiKuOuysiK/gzg2TCWG9CKRWY
EaGc5qv51QkEEf70JAKbUFFDYK9WS20bKrsA9VFYdtVwwpO9aMlaQK88ZBeDBl5R9ADmsx7NMmcI
fvRpvJqIbz0r6RrhDS0S4CR/58Zfnrm7IdX+ZcS4kF/pIDvN2S8rhbnDRMdRPuAx3YND9HbavmGg
QDG44v3VX1iLWnnEtJnQ5+7VkOjsByXgMv+Mhec6QtAaaqtiqvS87+RdaZPZsmx6kDmD9Mxd39LC
to+wq6pownY1pqBLsLZ8ybu1DAPYrp4/416Ledhjb7sYMVZuL1Jey7Jvli/cZf4by1moqGIShGR5
YX/T0plGJKbA/UmPY0Pf0MBhBzq8kxD/yV3vhtq30t1Ybi6ZIZD+0fl1tZJz+f35NJLipoylgmEE
YZEt0cytNOkBZ9P+ZT8WGecbD7PxlXbeBNH2ECM3zKV+6GwWpUbg6EVOb2ocfzgJh96DCt+HiAjR
CDF/2jGgy+yhCeHKbgWn10wbnkA8YdjeRAU9zmLTzSixdHF8v9BUOKc6dvQdhVOdLMkqZXNLjrrz
5KanRFef7oMm9Ax64qwtYWQIFsveXUmtJumqRd3hxxhx1IP47zsnr3Fk3WK0t3Gowy0Nju26/6cS
bq39cOUUiAUonR/uTda7xdprCKlzQDjZds+Hce7il1cw7u+ovb1NBzCAFsWQ/JGFm2kNj+XQGWfZ
eBI4m0cMWe21PFY4BOclxhR5/L+MpOCI8BnzyFuHkhg8QgKUqGIlV0ag7MP5L0lD5DvtoXW4icgu
8wXILFYcm+uDXzA6tqDL8bH2WHQfT1jrac6V7a0aLvsVbSTz7KQ9yQcG+qteFlp95Pqx4kOhmtqx
f2vCItvKDxLbc4lEQ6ZVwck7nQvI0xuxzs1jJcgUVrZmF7BIPfJa7ri+lwly2FNRqcipwp7xGPDJ
KrAt+wCYZekgveEZPQPIpFQyJvW1jfEFHklW7gvjsUB8nCTelmI92KN2JGZ0yeOlBpiuAl9hzXtJ
PKofrRSKl3iEc2rSnSn0AfAXyDjXYkXcDhmDnKSEePQvhkSFnCr/dmheTv9+p40MrK7lr3XJYDyP
/gl+Xwc/a/P1ofxuv1zutvB0wxheblKZ2NHx7oOVAmOVXuG8RJ6339RLtryf9hgAR7zYP8H2n3z9
/3p3Av/lKHSkwTjGFpg2byA8qJjqrWXpsh8Zww+c1x1ccAWS5H4ETLf3CbIHqCnllMhYbxFLtR9i
EXe/CBfEF6dxtzrZBTzacFaqLQfuyNOZp36YV2WGcHgUp9wVbxrYwcpmGTpyBmc2WkLH/Ebn3LEy
GIUZ0btQvm8TFWcYasRr9zAgnpDraTHdzueGZmhLUPvk7CMWVqJV+UuCV8x/yfhIm+GF+EZW6ds4
U4xa0yrdz/99yvAbWqjfgBCWua/CPjyBdHCMFUgk3Co08kpug2gIayHyC6yDtWeHXwLaFkRQ8OAW
p3B958UereGuHRCr/6kV6ZvkvZ8I+zHyIxGv0LfjZQXoeu8W/cx6/llqCWaumbxABuGN4DF91t5h
JC5ijxfV8qU6H0Ymxzhcsnb/+ihzuNNRC44LkP5gdq3IxhyGXb7+w9BKFPgjPqNGl81rxvRZYMzC
tdU4AYJ4bND7Npa+R6zSpSUD3ppk8r0lYJODlu3uuDErsfyzAbSCraG7quXqDH8e+vTogSgRY+dY
9JYE/YmnMgHGgwF4Gx5HneLgYEoklmnj1rI+yr+qhZu8aAKcxOnd0tocDJH8MnXBQVE3IrNOkE8r
t7A8gS9REiqL5BDyxoV9E5BIAtsz52btO3VRB3lrukodD566vnGodl0l3K+VbgZtrv49TKHQJ0Ex
8J2EOU++qyH4MdEl6BGxkDH6Ar2xZ0C+hNkN7r3jjDUiV6YEAL22w16Rhh7O4Xc2yLCwVFnh22vT
dnm4hcxO+Q0IAVc6Zn674xRtpnOdZ9BWuakaSGxKLj3XZf59rKMXkxDVxc8kE8KZBf9X5Juc2/W8
EojuN/NuqGaxwWv6/alIPqh9yobcmaohyzEjUzH6IBmMzAZpfIYhNt7PVh1qKzYsY0DFxnVsCw12
rElWyytc5JcYY0DLN/pByC0KNPNhmXRG+GytP0EU9eO0tzoA6hYaulxkxrEkfZzmYN02riml+RKd
gPdxqUrk4WDK8JmchzeeLx54Ugnslu6eZOcjtyg+Qh9S9KWGXqRPbzqyDXDlsRyEr2ZJ1N5uX1ce
eKlb1pXMW7V8H6c3j46H25azng94cASJZoYjGy/rCjYQSTDR3DHxLKLb+QoO0xsT23/LSGW6JMfi
aVgFwkX4Fg6/S10CkYZwZB2IqhE/DA/7eAqFMvA0WcBOAiYw//igCyvmEduj+DMcag9xa7yeW6tF
cB9kfA3isuG78Qi8dBBPh6I29n3bVgPVUxYM9pG3uqg+DPC7l6JMEHczZ0Ti6Pj8Lsm0l4xm7Bwr
r/Hb2RvSbOlJC6qqgf9ItbMRp3HE6ncmJal+Ggrw4adzMgckY8Qo5z4vEhzr8xM8pwUpkFotrxQS
yDNAOPVfgJj03CAgl+uYoMzl/lBcIXxp0q8edW509UDnLjNd5lB/3Y2PEB58Io5KJuoVbmKBrS2a
GK65fJB5VKRRkxj2EueLy1sHaSQRbCBpdQue32XDRxVmGT8royJ7XrsHVaFtE5fhWDxZBZgWn3Zt
xWLiU+gZAoO415OixCmXwvaK/xo0lTLCoJwPBwL/DW468ja+22hxL0niAR/P0sqA6SreE/Um9xnX
RssI3rpzDonJcuz6g/CbZz3MvDZ2/3/aXVC/mFxjab82OetdC0TfseRUXsIrkeSQi2QmyXqrAYw0
ZYGwtD2EmbGpEDgv+NxlOt6QIQHO0EWtsYJq3He9HCWPDDyfRAqDHFApkEdP3kfUu5bRMmbQJ8Jl
pB2ar3R0zm5xIGeA/5ApOy9BuPblSOOq0KvLkBkEbQTanZD//0GoE9agxaB1vsrnt5ZtlhH+vSZH
fVFPsETdlJt5hr9WDib0B7MV7l89CXSbqLPsVy9MOmGWRXNXg5q3glZ2rkcCN5TnQSqscPjoxIWZ
grZVkd6c7hqfCVcDEfqPJdffBzMor5DicI5Wv4I7L+FdAP8sgzsRc+MNMd0F9D3gGLR6s1Pm56Pp
VKyY5zpu5m2qn8pqHf2z7IBvAxSgN9Qdbt6HY3MrVG1NzkmIzTL2DSVLWda3oNx/Em8cNtFsJqHF
Fdg8rUzo9WEmuhI7jpE42/uzSLmoEBX8PELl0vmkRusosHhzHBAed+HLADqyfWbOtD8178HB1Lgt
dHH67YrQKrtXq9doOU0YQES094EjTxieQnKHXgbm+dbYzFlrsK3KKn6r7rE9JLAfP6SIFEwjrhgW
kBzSVQQa5++fcZFkSlqlAtxCLV6MoA6Daq66x8rJfWhMXzoFVMgUD2aE2+lKhJBlLgVF5bOyqBG/
NHB6YTuCHUxRW12ZdZ0l7UtqDKhPzqqr3NtTVLzJko0pVW62R/Am+mLZ46XfqZ16pdwvRb3Ek8x4
7XDd/3hJ8kV5fBpA8ddCAQVzkv3D9xLDzl+FnpbjJrDyFIiw95VQayxEcYf6lF4c+C5xJWyhX6Xh
1E7VR1neu6NJcFLWmRJBBH77bsX+reNiUX5bNjsp7451o3Mbr0keZFtrG3D2IehzUyNYKDdvfI8A
iKddCwD9ernNM56Nq8txRoCo7cDAawfMHYi5PnEb0/5G9g1OVp9XvOzZxl63HGiCcFuTqYZ9UtPs
rIR68dcdRAe4QOnC/aIdPjLTDeiyzz1euSaEA/WkcCC0AELguPDQh+O3+uQN3GiiDuBxzCKzUOPI
b4K9wkTZ48Zft3tTrKpze+IeLBRHSOFAc+ReLXavJ1F1jfdH2kezkbyAbmNwGgx98tJ1FrDxOif1
qeULXrCsGHk/oE+5e36jgkxgyxHy7Hc+g4gVSuGoVz2AdcN0i6susLPIYNC2nYBgGp5EAUpe8D9z
iIXQE6LllBqkOjMtcw3wb/ANkK7TuOXA8ulhkK0axkU/EJcTIA3XnKilI5fOm0/PV/bcQT6rocdW
0S+Mpu1MDJdoK33irl4it6xJNfe3jVL7TYfDDairo/pl1ab6km2uGOqvnaP0M1avyleiqbPduhi2
RTQ3iJq4dWJrs8caAyHe5DbtqDLzWaYPlGCjP12pKd2E6JiE6M/TjNDG7N/YMByM/h/16ZWiWxID
K59UEDFaXwWcYJos6agQa6OSzvW2WdqRy7Fo4STgtj+kmFHhhnN4BMM+U4o4QofO0snAMWhDYZNP
SOtYcnfbU5I+i+IWrLDEmo6rk+2wnKS2CdCEkBQ3ecfzsB08/b06o2DsHzlOz+9AKa0h6SsfXltm
A5TtP3Ul0T/foN/1yd858dZbOYGXdjVtgChXyo800UgnNFUaOSF2hc6INDkc46qAaZS1hxYdxhd9
Z5uMUOlOD+Rq7poOHwBY/udXLG9S2z/3aONM8KISR9V2Ppgqp+rSCh4ziQuaBEGM3yTpH8RmDsA8
VrET9nidPMiHWDgMrW/gRiB+/ytL8n+33YhVo1eb4tvsjICiuKzMK2uPrausis/A4pcr4iSLIDh+
bFarfUyDXeOKueZ1Vy3+p0tUjkXYYw7MCXbIYvUVX7hR5vx/rfU28pMMyaOs4Zw64qeQH9c3vLCY
9l7pScprVrK/nZc+CLVedSpI9mMa2takjJGERx0ObQsrHbMdwhZSlbKXtt8v+kJ20It/U2M7lMy1
6gWhX4Z7vWaChtzaIONnbxRWoFmCnQoFgDB8VBHR/H1er7HjFxtSee4PZjRqxuU/kJ3T4c/r+gzq
p4qZxBVjHpUAriw9gKz1uizfVr2Geghp3KbQcDjnOelcqZjfGXa/i2bN8lkFndWRba/LTLrHtGUd
SdBRu8lPQKUlAT5G/s7bl4b3Qpjm3eDHRk9wNkMf6OLvl8mL2V3Upq/iZAKL0j1+lAFE+0TPlknd
lW0HilE6D6VmvXEad4bGGG5PIioOQc3XuojV2Ku3sEJLcrBsteW+LllNKQeVEi4wMsDTL9uhfXXY
R3gto/LQvywXojHRTQyWzk5e4liH5Wq8yZsLm9ku8mIjr4Tl696FVpJcfGk9mM7wcwnUipbswDlu
EAd4PLUAKgV0H4O/kk0vqdNOMZr6vXnQQR6eJtxmeredAu6jUdBHJHBMDMAWHq5NlMwgKkcDX+U/
Po3jAj2w5sl+5R97MUVbrGCqJnSvW6rxfoA/ganaNV5/bowcjkBfiruwUbxAusFS8kGHPVPT3frg
5If5LXueFoSFUqUrlKuBSHIWLI8ubmsNENmwrI7W4AfhcYeL4gPTDrIhfy5QplrGj33ff6YveMIx
knYSICmd/xuP+b28d7Q6H4h+qel8R57WtM0n+99h55qo1z5b27cHww+KceXm8ZC7CJ56sWpLQ+Pt
qopWqI5bsyDsvHklrOi4XtKPBwfS4GZp2R8wwczOj2BAZ/x587ExRIBXaZYkyeDb0xjgJ5kOrqa1
q+AeRL5I6R0BFlpyIAQuJtflcVYm094OavduiTQ9A0izhjUWs3KgwRldxkGaHDIv6xWMsehzlruX
4L/im30XBwHUijzhqVRc7rHReZ8F2SjjZet8tc40KQx9ouaFrmoRwJIc3HAP60g0EaOoJAH6obff
0TdM9OEET7IpP639fswHk49100Hw0H4TVXkacO3vwcxm2dnHRDPNHl65duCRVuh5YXpLth7ZQyUE
pxMwuob/pa82oESA1pHcJMZxZ7T2ZSFlZY4IXEm8PfkpGj+ux0XNoUasLgn5RxiLR9oWWCmOf2xa
4FTjOltA0e82RDelLh9Jo17Uzo0SGxkijudkZdd5R+ANm1rufOQWzAlbWuNMkkZWxJ/ZuIOpWJWy
VqVplcUtC9nPQNslP1Mz+vE6TAWXOEOQcJpSHT1lAplCTHCsp6SHW9BtYxPkPsD26VwtoFkcQMak
M/1N/5ExcV3MAa+zYouGvfWGnYrX9LwhpBl794az1lsWxLN7RUPsBj9mxzeA83bXbxov7zXOGdkZ
7Gww3ePe9FprR1aR9kxAH9hWFpM5/Y57zYiVZ16s/etVleA45/R08JcU6eeZ0Jp+T73X19+5UUm5
NvrzXUYN5U31X3Twnfmwaly6it8X6okm6ExzJ24lxufrRV06FVvwv7wpUhYE5OdkGydt2ZgrAQBZ
o6RWFHooNMLosBv1RpeMkxccKkU3pWUoWueR7p7ADqnLqu+Bfy1jDE6X3+KZBH+sEC/7SEtul/ZC
QdgLhI3dq8rkLzhtwO1Ao/8bFR6LqvxAjicqzN5aULjEZPvT21zuNnilznulHZe90qAKJTX4Mj63
dkyzkd9eVdeDcPopPZR0fOAWB+bWl6DwcSuB3rvL4L6UR9N6cxZ9FhyzOY2Yt/CsFe9pHxomBht4
DMBk7QwXawy75jSQM1sUmJP1j1Sw/4E7oHQni51LEvSiHdiBiohKYD5ZhhSpZp46hHBCMyWFmxqV
MF9yR+KpcA9vuNCU4lkr75e2ELrROMGdoQF5sQY4tNuRGo5PELjvwvnfaLn5pxXYME257iucqePG
Vc/LcrRyWaQMcSj6rLkJ4UIhL8r8OXuQotKcI9UkPXtiQwxyEhrJdXU3DN+Y2XXn9Pu2h0/GdD+x
+47SKjEWzCeWTX1uzWXlfR7ZgOCAitG7U2xSihpqBvEwz84RQ0QZjhWpAQsvgMFsaDcD7+ADVeBh
CRk2l5+Xvg+2YBiRrLYitCm9qjprY52JYjFYTv62afLryExeWa+0o+NRfCOCx6glI6iwSAqann/0
R03dTdV5APDUhPD7hwJcIKPZMgRqxHomqa/AmimtgwaChiWitVkrhktnyMppMiUAI/G7hiGSM0qw
KitdeXs4Edj7mKq4qZVdx2v9Z6J0XmRAzpK3PAQ7t0BdaD0wWG6oAQMJjXM2jVNQcE9Q+EN8W2Lc
xJFiwYnCa85fqfnH+ebdKPUNPbvM3IhogSochchOCKmAzZ0PbKnCieSlPdjkHfTjwY+9oguWsxZu
XU780pK+Xg5Mc/Kq5ADDzXHVRLIDwvaCh/eP8wVOwTeMNAGrdCBgnOnOOoHuEnygiv5oP9IrEGS+
nRyK4AhZPzbVhD4jr0UH5u6fHstFqJBf4B5PNt9JtfXHBcn2ChpXB6AKgC9ZRuW7xIOXQmjPXvIB
VT2G2T5SbOJHMZ/uenZNwpq8d/8aIEpHudLCoP17XSvdY7Whsg6TXbEMbFQaWwbYwUFPTj7iaWGo
24WTzBCH7t09B7iLwLIgHFfgVigqH9cu2Nf35BkmdNrNzBiJvFRec3r4v25UQU4MHH1LBdMhEEKz
JP8qF47KNdGuHp5isbsASaCkyv8krVkL+tT5Op2ffJCdPIvX8BcgjV1pLatvu3ids2Q6wALayCU5
iMZ68WD12AmHsw4w96sOTOjxkdiEzG5Kc50yjXuZa9grkbw6MbO7pbWGl6NIPIJUWL98Hnpg/XBG
uZTX/fN2r8MVmsgkJ5lQ5vX4tPf1F/KIWJmMSrCAXQiwwhppeTU8lBqAI4JAVlmxbpYGLaTmk6sL
+2m7yYWDHo9AIdQM07R3HpOa/BZ0WbpGXievLuPH+AE90Pyjh81NfQEVqwgPmF+m6JQgQ6+RE8BM
fev2XTHwxvwxzvRapPetEvfT4QroMHDvt9x/H7AnOrzAKZk0UQnNXXA9iFpaP0SLBROMOHIPF5sJ
LY6jtw1g4U74WcyYbP2FKJ91CXLVMc/hoGUrhTzjEJV0JSqaVPM5PrXlSdjbtSNyA23OILq19lDk
LClUOXcNsMX8Nw+fUE90f0FyzKeGqtFQrJgeMyT/BFpaI5/b3eY9DLPEyxvTfQ3lct36+ymMHkFu
YG0WSA9WqrjIX2N4xOoZQBZVbbi5DCDpGOL9kNOBMqLvLiqi8DryxZzepKymCguupxTcLye2r8bk
JWuGx0vgdYSmFhsOMVZwmAU59lGbxHDIFxsfc8FWZZpxz4evtnfMYBumn0ODKyxi5WV5xFI8IkRP
OCC+hjFSGhG2d2O18N/2W8r/i/NIvj8iWv6MSy7nO2WZBnK/GKY0cmnUgXtBRIUcWn18GeLm2omv
2Z15CpbtUFo8SPjBt6irMINf9cDg5QV9seK37Y1HOnTOhSk5//eUbfrRPklbJ2DfIX/w26R/IL4F
UI//26UHLtjG+vN0wZqDn/l8yyAHuvFt8nbGhSiSoPmC9ncRvB88Q9CrKKkGfimMldmWpb87wr86
ZphYGf65kWp8uJruc1Tba1p/XVCS+unPGESHPcgHf7ojJ41zj7QOK6kh0W0UrrD21hrMQ8jHaxyl
cme7qDQ8bCNi4JMHSxAuYb0+YRsXvKPuxgEHQTrUXavsW1bdZrsOEWU6lpnVh8eICKQguiwZnUSm
K0cy/AMKZZbDAVqghI+CNuyfgNy2u8BdG4BGo0Hd2Ctr1BGQPMD2sL5CYjH5bzyeFxRtF9dh1/zx
k2EpDnXBXDG2mlfb+fv6PL/ISFv4Qb0PHTOFBmERCuL7f8mdbMINjrMrLqztN+6PTTgtv+/uLqRk
MGr7pVS0dGUkd/ruQYv+frQgI4+8W4buXAOx6/tK3mrBVngHdTxR9kWaPP03n2Wj2RS+gBEGhNou
k+daSwtmyN9bimAMWkiAZVFnWv2B4ZQHrKFc+S94gVh+UcUfe2Y+MaFNooC1QhyW391RsORYYbM4
qpKzPl8w9cFQW5yHiHF5tMLJcBU0cvULVUpG4cGKttMTWt7Mtsx+kclwdkW8/1oV5XWgEvfSKxV0
kpyljv3/lgi1Y5E4jpGQXBYHFvAY6KmwKEM6DSA9wspsQU7BQRTrZ/5KizAo+lbDQaW1NVqKbWmF
BzVb/9fTI8o/fDy3dPqdYMh+Qd4k25hPXVDMC6RJNO7kXSfxHakur5jj0QD8ZwR89Hi/92bCill2
oONgZWuyQJuWasSzGMQ2jSAWvGTR7h9o4DnO58sjkCVaYgEJjxkE0H93/ClNfq3VLJ7WcEXB5wBS
3Pr4RIxtVkq7sWDplDY4/0meNfWrGTEUEML6DyLyzOEdwAIqdrb/poEYP0RZpT5FFlDsmiFoMLmw
ZOnaq57aAWbFXMwWPM4ek5Exe68H4xKCorM3o5vPN7+KDsrIo+a9+XzuIVv5AUvmyDf+1cdASSd9
r7rMp+hePJElKlvzt7y/9O5zlg8RiOQolo7gJRs8OEElKG8RHNRJlNvwGnaN0AlcEsW0Q+iAf+Wt
yr+FD5OT1S7KsSnzFKB5Vk3WmPNYZKjmohHmyY+5U2pml9Ro+g5zWMkmKRF27F5Nez2Zge5twyYv
7yJERLv+8X6dTL/qtxqJ75G+HhF/aUsBnIf3AUbKemPObHVtfNaVpx5iXYnrn6+bzOpDiXUcbBFz
+2MItz1/QGqtsGS8EULzEcK5LfFOafQkUEnCDa8p/TrM0u8lIsJLmA9STkg1wmG8S2iV2qETr5YV
g+iVA1oSvGQ/U79GHo/CVGo7nUA+nLtPr+x+i0m9dO9IMkVt8CX+ur2TWSlDeYj7n4m8tVbifD5l
pald8rL0DKWbAoP/Pz7w0/0G4QMMZztLjTLNVWXO2HKPACc6pF0ZVvp+8kqIWXjb6MzTLXZjVYx1
PZ3FldaItoLit9JJ6snKSvUUmeDgK4xK7R/Hj+FcY6nGSLK47uz9vrW0KEkZpPYcfhIL4zr/epx0
u4KP9b5L2v5/aqQ6G4MGt3B2CN4NV25l4D6+O/5aXy8qCtEnY4JmPKkZfC2UejlWBCEXMTYdQSUC
CsrDDVFVS06t5VE89yCOZKQwwVh21sG44Q3TgRIUSCpapW+SgGPHgNI7T66XtIrj6FlEYLHNBGbw
5hFT89R8+0W9pis+1x9974I9IsDwoG658PRNlItc/We8yW+RFHqVgShCNIKcpLk9yuD3LVB8Obbf
bjSycKQx+dGs7yGQxUjfzJQuVl5taczXGs4HV/TN/m1wtc9xyBXHIXs7a3OV2L7xPnQiexfAE0uH
L0mQ4cZ3099Zo1VKJbJEpz2KnKnv7J/Yf+wlA3V+jgrnnqnRbaaCmlENjJrCO97FfuQFz/f8kpME
X1f5vEPdDGdORhuWXBy3X71UMNKpQfyxgSV/F39nfoEgoDjf99NrD+Zbg53Emqj+UnbJEWf0mAw7
u439M0nW3GadnIehp6ouyqfm6K3GUwwijq0x1kSnDh8PZuRYxSo5b5VEgeURkgWbcAtp04w1dooW
5pbzEM3hAzmGZNRVHOUl7P+IljGlA0OxDZx6CW/8dy8ZWKSOlQF/n1jX1DMvNc7JlqS1JDWdYkXS
37BwOdms3XlxwMR/xlfgo6eC7gL1EowNAEizPY47tcRZpYtwzVEEeGInczncuWhvqqHGutf7ioHQ
fJLMh5dVjeDoAa+4pb4YfTvBi09IsU2Y/P+vbETzU2JJHlgK+mKGUY6OVtWbvjUxXM2My9N13E+s
TXNDY4EhpUYER0XaUPiUnmbhVsGkM5bNavwgbh5vfdXuMyotx/qeGf8QNzqoEFQsqa+Dp1ThWd3A
1NN8uuIuvGAEFaDVqN++ypIE3eFRZMCwr2bQUmvKJG4o8nAdAu7Ll9RK2vv7gQGEiR+8H3NgLvPv
pFLnZAjw+CGBXolEBBvqTmwqhgWmGc1djTKYJf5zLvV2WKUbh4VpG/PMqxbmD/lQMj426XP+5KVR
ZdAbzEcRBkrFrWpJg9z1uF2fyD2DPnJpNxkJfqYNmgUVQ52dwU60L97mCjE/8zjFS6jDuK7rbszJ
NufODbkgivH/L5DFRkoaoCKEvahgB909nuSXPNza6Ql7GLlAV0GncpjXnVeKuNkhBiwbQ5aOaQ15
09uKaHJnX85pb2i77g+ayFgBFJ6Pc7P8B5Eg6C+cD13cg4ejn0LwN/h6nQunq6Sbfc1E4xN8LzOF
NQd/KBlUcPh8aPHYs5TDuRvu9m8/OvsdA6pctlYBK0BthfTlJC+Ic4N/EUxIFVnyTGWY25IHHgS/
9efUnbWjklXh6rPyj8Tt1KV1qpgngknEyh2mvXA3RPNh2xOg90XgWaPDrONCIETBdzB7gPafO5FH
MpxU3pfRSpAkXDaqMrHnbLubJQihhYS9cPpnsXR7HhUPdIt0N1cmHrj8O3YysxmnIRVZ8+zUHVlY
yjGU5QPECCSDFMUZdvm/ZIFggaWO9N5GHV5JEsgsLvQ3Jd9jdZXVQxpD0dU7i+83L8/sojUPJ/Oj
Wejr/xIynXK2FM7r9xQgIXl6pNCXaZMciZ8wfJh02JdcW8lH8+QHndcYaeo7fcDZHfvXrRWIgijF
ml3reek3BCVkpfaaTtx/gueqcIPy9m8dZBom9ZrNOYCUaT3/VYoRfPp9+1VT0Yida8FUauZqbhUq
MOIS/IFkhiTjTV0mpRBj7tAZfD73U86ijhkVYeMBHua+LQrsR0rjxnLmkhoSX+tszer8qLFx7hkT
jWA5c4eL1ce6Dez63mHyVmoJew2BO3NA21ty2Gs/siV1kLZY7duWdmI1zcjd5WrtldTkeJ/TAkgl
TDgUrRHmZJ4qF7UDQ67/J5k7NnnzCwRsBxgoIoMyT0cX6lLcPf5pgVMyVFvYBVIf52pmWV+l+jqb
bC7n4p/x3OSB7D+DKSfUhILEm1tCzKZvCpsH/zdH7exX8P0dqedvMXigGBZd6JGn1WixzBBVHpOb
+LWwSa5a4BH0LVOnwwX5NIioERfpfynFvyhVykrxrrZArOMdhluuP4sBv5OEkwC/pJNvW3WEeICb
vxN/8E2XZd9pM0emMk+4Rxb6DyJ5r4RyPj2+7itd8wdnn8CIMUjbzOMs3BR+TbcjPJoXQm/uBpYr
pmRqD5zpPkQA4fL4o8flAO/ok0oxVTxPf9iER0uBAB8RC3VXwGu+UIUMXtyH4sNyWxRHKc/hcr8s
Mb+GMxBzY7LfNQILcMbxVyX0cdY+lcpY6c80sX9Of9ma18dR8tHMYSXlJ2bWFskUdT6U1ErHQ/El
06nTc/9RM6n11dzSbhFSc4RYoUc5MXYW7hVfUG/abYfBoHRQufxanCaka+5GukOXur4JnjR80CL7
kIwR/h5htqbriv2PIamIFRdNmMHAgJVclYfSI/iGdttXbH/bp6SdDgTnAn4WgLsTcg1EbuvsodXf
BuDZ7u7mQdOTwAWx1BP+B6UIeKzfzHLjgW8qpznc6DkeC9vt9IqDuJqZgAjIlt5f6SglhH19XVgt
BAHat1pf6M5LibLP6eybjclCOMwAAHbKTSIBu0CcJ8qXL/XeONIG823Xs0456qp1OaMq9p7bQfzG
+gXAHv40NFj/P7RgZGh7ruEAJ0O8BD8uKYdX2TMtAT2nuWQxH19wFH5/vsdpRKFn/QdnocIib5B8
Xe5VGaVbc36SxNc/eVfWdg6v7fG6qnQzLjEXJNbIQ3P37mZuOzGtBIV4oTGFVhlW/tHIIICyXM9A
g3Uj+5X2iC62siH+/LUIfxnxSeySzf/Kql642pRSNJiBYGOYUF0b0GeehXJ0PtOPPnqvg3hpl0dn
1F3k9BKf5e+nDIfgHEHXO+NA1ttIPWLpRRXcrliJnXSSnfdwEeVpir3EjpF7cIC1qQ32fQKtt7Jk
StYgD42xNiQE7jUBknQJVwjMvsg6Pzl4jsFVDMBP7dE45sMpmXDw8NbiLih8MkbrJ/EIAN63/H8c
y9cAqU0zHkJy1rrXrLxigrm2ZivvGYU+njO7rsp8qovS67DmjHMNuH6UI0THTpI7tbYjpclutCWi
eAVOqW6if0Tq0IaDVaZruOOC5yrVNrhIngLOg7lc5FtA2Jc/pU370TgtDSXazc6VHuRh0Xm7HMia
/XQE1aWxtIlR4iWuecZx6bnP4zcGls0dMP7i1C2GvjmsuivMjQ8NRRXn2AX6Mk4Uwl2QFvEZoPnS
XxCIkSanIzJYU3WdPkQsL4tEQVJJ5Asy3vAD4U0n2qCdBB+iaibd1UrSwFGMa4RAIzyO/SFx7CV1
Lk+qun+PWB7Be1PajpRfC+s6aLExQv+z5Cq1CbWoRMY/1zvBHeL4jqaoJ/yHlWkcVTSBHhkTNZhB
IqMmHv5Q+sNC1uR2Wjg5MlZfwnrlKx5RE03ViPa0uibsyVRxl/UH9Zpnum19MAAa+Fq/1CtY9iKg
sgcrlrqk/BTUXL5HE06+IAs7nud9GoENmC7Rj7x1uFfKNjaR2cscUQt+zjNAgGgjsWhsfvwE+itI
mZxLDWvtW7LKGXPXnWzDQd1xI3xhlFZq8FLj0bw+gkuhvREb3vCJyneM2ih0pKoIqhyGIVkcG826
kN9MDrLlhQ8tuBVNtF+6OP75KXJB+3nUA0Uin1UtXSvB/2C0MjJ4vghXkXfAAdQ+gpVdy7SdSY/V
e4KpBQsKsVsyx1XowwQ7svNdVlXx55cOWod75kCqm/ip6I6SZYOBNtIq8psHB8qDKZQ7YIZ9h/3b
vqz6nzvt9Jlf4O7cDA4LSsX055qx33ovZFhtmSjg8oWdhrImsuIMPXYatW89FeuFIsYIR7WFaZfA
cl+yp2FNOr4Ox/TuteRtAysVrFrHxUr5tilbDISF9iakelo4jweGoHffJ6hnCEjcxIE5bU97wlhI
gJ1h64xinbPeIegrQgQefksbgdTsPxHug/nHNUopy+e8FBHQIvJo8N7RJEmwFBpRozCLzF4pnZhb
kWyeQ2/otpS0UNPLtaBSU14PVWL+xchT+BRFvUNoJs75PPBTyxcBa1xaRseFp2tAQmK8Ir1k0KjK
6Ml7NOM1tSbXIyoop05uLOnfVbdilBSZKNHyOmgGCKTcpZ439vDZxpgMgA9R9KZociC6NVG5WJvz
mIgGAsTWhWofLvCPiOoUvjKUBdpB5bYq+rpedvYSFgpAytMtkogGemZmNlD3NIUwzYMBltpCFwTY
p7BZbGcZIWdhcBSCt+jKjiqHklvoEgnCFUdTgsRBbXaTYyon8XKxio7d7DF6B9+io5R2oPR/TQ27
coJNw0KktL27RjATNTobFqDgBUmieFdUjzPMmgcKW4hG7i51Cl63qluMUIg8Lk26N+/pmwKNCsMo
g4T1C67JECVG8LDAyfU9eiVFViR1IzUa1x64MG8ACBCZxLgw35rqzXkwQOHDT8Hvt6WxoZqsXeGc
ZHlAYfqTyiItWnYJeUX5oJONP6jHnuMjjU3TSMA5MJu20WZVPWjk/sjS5idacoaCxdbCXUniabRw
E+1T+/3E3HKBuqGgmY6lqHfhlsRszmgHNwV1UN/MBnbZKHGU181k6yRPLMncZl4Dyh5XPgJMsusj
5AcFadmcjWrcu+mhq2bYV0bHUye1rpreTvQxxiGCT+RE1pVDG2uHmRwuRXsL2tfHYtd3gU39m7NS
eCk0AdvO4nQaW4NMzjEWNJ8h7D/0j1GU0kBEp1ANIOy/XE1z5dDBRfODl4uwShW9NN0cuYO/feQZ
ZvvkgpL6Flh5j1Ofm4V44XAnfyKpGdELdifxesIfihOxKsCuqBd9eTkLg/74hYQxtqBXZU2cfYCb
IrAkbDM9KNinGnT9drIVP/UGCT3DmhgFq4civVQlHsVZrZPIz0NvMQcjWP6QULw5CA4eoYk6eiM5
EuuEqqIGn9oMR9MGulS++MJ4ROJaUakP6PewjSiNlcSKEBjplwnPNLAHsRBQcQDkZ0wZzDoumUbH
5eltmK46l0Fim8+DzT0bMYyIYb/UBQF7sukAMdOY6y0v99MVAcIziMIw2JjhqpOuSP50+vNSROJG
HsJK+hHkSh19aWFvgfBV7qtHkqdy2OirF4agPceobYRTEm2LUxrAY2jp9moA+465YmEcplcdjTfO
szGcZlUfrjZnY5i0NeXTe31vDYHFoEk4Pbi/OHHsRHG08YJdv0jZ+PjRDmHMII5PIMPVdrXtlpZO
1pKzCBcIB+f1QNw3DAMKpcB9MzQ8HTXMRQ0Rqmo2k3uwqlECxrEgLH2RR2ez3zi/JtyeyWFCciQ/
SXvQK0XGPviYiR1+e6oOWmi8Dm5cdbwrBNW3gQQRv1M82zMxul15UsjbIEzqNPAP/gwMwrQCr/AJ
mAD9lzv+9VbkSEizcfa0INB1WGk8fxkOu+IJiyRdKTWkmw1Y3m1KGgprL9Lb/aSau1HknGkEpnt/
1DgnsVJt2gkgGsoXwexYMrRqvJVJIwST2CCHIqZuCr5KBlw8EQdfQvy+/kESOj1w2InlTTqtwybn
RMGS5LLMCI4L8KPLAtfZ/q3/1K/+Os8NM1/6iPP3vH1/fxqQfiWOLJKqMFaEOte5pA/crMrufif2
tYr/x2TDaSbH7oySHlAAZubI3EPycexqfPeZMq5rfRGBloyZHRGikd6xkcgnww3HyQx9c0k6v4ON
pX+z35gc7XVZNmiECIAZAFCLwxi4K3HVVVBg3jKXqn2kzNkTjrU8RqH/AZbX4/6jt+aquvqJoYks
ZKhBJj4iYlZY2AaPiWcgJvbP8mfzykufPm1nyVEH01dUAlAscHdbkHHKzuZMsoauXluwRaaat3mG
MlKmh6Sl7d0NgWLN9oc4PuVF/vhUHeFhHhj7VjhJVfxogL/dWVAjESc0X6mfwaawOAnpCKZLiy6C
xZgGtalF4qtoO5v/SCkPp7iw8aFM+iCEBnKYlvG/5fBzqZLpvBeNO8Xoubljb/3MWOpC67Kw1yck
XLjJEDphUQmvP4euDSqBDk69S3EZKb1I5lcE6CNRQ/y9OzqKbETZ+eXWBpRkOayX9DlOc+4o+qyS
0VFxw3j/ZZTuAItsBXj914fg0XVNX66SlJCkGOp7OkOpLx+6FDBfyujFROo2UHTL/hz3zsbY0ycP
+D3AQFivNoWFRGbaUGIQHBuA/OpZ9z5lY+a+yQSHOsqc3K9Qkl0S9WLoBtDYFmdKmy0ROsVUv357
1zrWamDcCPvwLnJ3INfr9zBsogho5gPYgq56eIClJhwu7Vr9jJ8P9kr0UiaIIK0MG5AxYqGeFKtd
QZXcqwQmNnCKqZWLqome0jK64MKVCNjy2vp7oiHhlc03z8HNgiXCaudPpeOf5W5RsNBggZVIe6WP
E0XSpdv/0Hd1DuZTdGNorYyvudsS8EwoewnCKFKCp8pg+QI91wQIiFmHI4s9mYzq3mG7FNxDGAUr
qKoO10GGUOJwO5jUX0RgrTvx9x2GG1YQ3P5n65d6orAXbSdZcvJrOW1c4P2M0w4vOW1zzUVffV24
qUDUhoJ6SlKtx8vINL8S5EvNDWs7LqWa/ZnrtR2P0ZjUpnp6x1DnBFkMzvEClt3ZYQHgURxCEpjB
/CLixlpoCbaEJJl2ONoxd2/VXemQszLhOXuVLFYQygKLyNsR2e1uHPeP2Seq7x0jrmDQ5bq47iop
2qAVwYZjv3VjxSeb5OimSUkUTbUB/09lBeJ3z3CuauoHwjXSI4uZAEB1vzkIfJz9YQsGFKcBAd9G
Cgj58On7NBgflNdUtrKRFEQ1qIvmHtlZbwyoDJa6V4iejbQeWrDjtAXMFA5od8cgRMoKAtPQ72zW
ekRcIkj8NwyjEyyrqSG8OkkiqufE+rcjMcs5CJqWWVCxergTI99CZvPFp4tnxU9nQie/aqJEUzRk
2Guz/EWk4zpy3xspBGUyepKgj2HGQc7B3Syk+mhgOLpHSiS753eJsQNPfGoL8Es7KZllAvK1p92m
U9DusoNj9YH4HbS/+kaMiIZsSoxy+W8pKnYygmM54DxOeoAy53ZvKBEhhA/Y519N6QYuxJpu1mqj
Fd3R2fseat4e/fDEyEEVlOKQOLlEbUdn/5CSmUE+9FtP9UHfS0lc3TKKpKbOov9NsNqfPW0EhTR2
NjjLFXe0mJxn+tEIItVLp95hDd6mruZmHkyTNXOgZAl1KgvMPC4O3dCPJwzilD62C5alxaUjQg5u
vKPHyaZrT2B5zTqusIm21d3BiDP1x661IfuyHAtn3JikuTgOvXm2vyiFtnqVPvZs9RUZWIyEoMdT
G9xMdKIeiMfrroGqE29vSIDniOFRRDDOBFBqj+QD/Co5bXEHN6Iepn6PXmxn2b5Wd2UpGkSh8bcR
mfx8sK4YHPrkBf+8SRhWj8ky9athhU79ZjZE8ujvqJAJlEZNXbaQLv1cDhGMs6fWUQQM6ZhMUKB2
pASuHBdHK2Z/3xrZTQdd1DubGOWPfsGDKquUQXA5KV3JirSJVgADE5XyEspyFIlOZBlDM0h2ZrQd
6ZKBEkcemtVo7MNRG+jOeWcgjLrkVoGY/YUj9vH37VBYhvXiJVRX2CNjptb+bW5N9WqF4t3eQT2U
zY1ORPaqLd2YL15R9OYeQCrXkyDzK5Qtyqx29bqkRlCcfTo14D/fjJwjomDmlQxt71EQHyA8pLu1
+fg8kBZ+t90VDOoPTBTgqEuJx1SyKhpmKtJ6ccgET9hb09Obvr7xw3iGmY2MHO11q3wLmOp2HUEF
8Fxl9dQvMLceuqDf4ZoSngbCk6DoQrVD3+2GTB+LZ6vxGiwnyPqmJGKaH2lW/fIvLzGfpFdZjby5
fGxF0LucDX3pQ4ocyLJY4gQ6OynW9cns8Px6Tsy11hCPU6+EweVNQVavUVENIVx1vRKR8HenmeQs
HbP+VlELoSmhqKvxpHPaPELi27EuAxNgGXlzQUNv952wHQSdYAbmPXeGzxGZtFQ4CD2ztgMHUzGY
VC8/XqCwee82mCOox2RCsiPSIaxMKQCfIM0hlYufdhDWOFz6j22txrIQqbfSEXYpNuZyyB+QyHan
lbl1afrLU3jL+Zbt+ndoeTyvx0HCIM66vLeH844R9JkHYN/BkMaQkXYj/ro02IX+cDrQ3x3nFcEz
cdNXabr1E6KbNZrpwWZQ97VbhMWKgs3g7Ic5t11obl4WKjw7NAhkX5aRluhGf/dww1Z2xRc9NCcm
zF/yVuHYoPfs9QM+Ml+rArmWcBq8O9elBhPeU3vwuYRFohavGHajlI7SAVmjdr2uowsfzlU+zUPK
GQnEJyQ0tjjpLjR/YK0BSogTUNCMuOs4HqVQhKVPNEvQ7KFQeB1STjpxOxbBy1fkJEMwVlEKzBR3
HFE4uwKl2w7TTByXoVmONSv3mRCD2suvwvv/xPvVgnHnYMEwu/eRQmEkLdZFLIzJv7iLJ7JxT60e
+dXstscEmR1ae7GxphzAzKyntjfkemUGe3htP/bfP9i6TnwIPiSUugMmSi4ZbkUlU/dKrFKVLEuK
MhGFzmqfzb/a6MY/df5dRXthtELSh0STHXQw6Fjae3Urb24C2f9uvJ+e54GrPF/9X5TljUBohlaH
lAWNWLSiUmlRG6WWSOO8rEhCqCz4WfWYuimC2fbltxtVfGjor3N9+wfFkZpkoLXTx93HhliaS14T
Aa0iWbO/+zCIYWabjZuQ5h+izdIxs2X8t7aYdJKvnVa8ss0Hz19FYNjcnsq+drlfSIJiF4i3r87+
Kjc6v5gBhyl5/IyS774u/iM8KQ+MxDifdQKe/+hcYspCtAPzrj9Wq8hGpp6K0bD0sHkvs1URhR6A
D1ulsW5vniQYfMTe2KHWCX3KCkbek1HjvP7mjJCEW2LIKw4HbBOC2ow+lgxoEJb/eic1HgDmscCj
4CDgPdA0KFvxc4JkCj5zTqkzmrw3/KNHPs+1JqK6EWN1tEdH2/cCxh16EmS3/51JjktDoiX/S16h
gh7/5qLDr5JOCfSsHipr4SOyWA8DWEVfDpHbmc021/Kop+zIjJSC9VVLfPWdMSGCYDLanPS6K2CO
07LRq/6r5QHVGWfIkmdJp75A1HpPzi0axuwHHEmwsktWwaTQChohu67ELECO2dUMBEc09O7dFflu
xXTp0xJUgjkXdR1ogI8XWMr0QJTzaglMwACkRfov75PkRcq8AR8+wIVYJGHnCWAto8xa9IvcRty6
c4atEvP8RgsE4sQeK52py6kbZQ+w1jy0LPT9pk+yhODDzDgaLkA4XUHjFo6VycNU6mHey9ArplCD
zWaTg2FhFliYabltHSl0ZJvDlkkmS59IZ6eXpeDkOEnvDPg6+lgmiKBQ5klnMBpOXjYoG8USm2WS
QNnh7MipIWwQIgKzhTeeH8ou7tjncKJL4d7x3AJG7kF9tbiqjIHnmu7/tBFx29ZZ4c3lO2r+eaaz
IzeDLvBgPgIgSDtIkz2jQ/e9YUPnTIyEmhKn+3+A0YCIm5ewZMWomRf/TVWDW0LVpsdKiBadM4G4
KuYrmbt6Ehb7KNpQpdEGfzQD7f6B5gGOeN+GyJAnyjwdMA5hp9r6FoM0n18yPgCokmLt7iriDFVy
AqKJ2XzFIHbJaBR1iweLtS28mnN1LqR1yUSrAnf1nfqJBoCqr+R4fkfqaPla32+lispVo3xuMnpS
gXuWMkRJXmuSudVBB4/9iNSV+i+ZK9PWyYop58tao/I/OhheH2z0KQ3KGN7OZC8lhHX6MuKWYWTV
M4/Ghn1up5IHCK/ERsAVEo8aUFYU9ul6+cq5CgWhblCBZwk2PNTPSAEpHVchCMELWIIjSD4OoJMV
yZbIQq9YSwo5D8S3JMiFtACVIxxSOh3x97/KvYM+O8VlxUX8WQZ5sn0Jg2+tGUYg8uv/ZbHYI4C4
VtQHuuzADvrdL6X0OhqD02Lumxs2h7J9kZ/dAnAHEcgq9zFzSxbps2vz1mH3mTE9W/nqqVmiwBZr
wNuqj6af79wNgPQAC52zI7zPZtNED1I5H5/vI2qx5AH+uQHw7VIgkF7jYoifZ27CsTMzbfe3kfpS
udMlZS40oUJ2B4AkCKAh+/9rdvb6pv7lRpnjk9UtndhA4MJzAUxhns6w2MSnwM05yF7dglF3OyfO
SKQ3s4e1poATyiRSK1u5Z6ZAq7Sxy3mOaOB3RaopaOuVImv3PBP8QtaiOFyB40M+U1RQHpvkFpg/
BeJ9z/Zf1ic8xNQcKbfbgVdnoUZc8dE6iXIi07mQarznXmcI/FZ1K6GXS0WafPbRsZKGMlq2rzts
gij+aXUjL/hcrt/k5JaCvl6jqPQCdOZSNpNODqd1K6r7ok1GqkgdhTASz4m7VgIa7CF7yHAEf4zN
6UcRl8kX3yWE6rf5PNQhU4hjOW7XNez3iEN0GZs04LPPUjF0LuCJNedGrMkUgydZdMt0An5BhdEb
j1E4GE2C4ojG5ApNNZiIscgGtkZ3E+DiBC7g7cFxdiceQf5wZfZmp+a8juqHRzDQVHspP9HlVNWc
QIRajiQ4Zjjn4T6/G6MfSynYGqPNKEcYAi00KRg04lLfS7bPgXHvhHuopIIJzeW+JRlEqnPfkAtf
dFzjn6BZz4UyiH1PC3dGQ3PNoDq8eUrrMppxkiLk9kbwDg1Gt+R8QOsSKMUXWTaFASPi6xFbQO4o
DnOKkkEpCdRDarAiQRsKOwWRf+qU4ghim6AGXQqMxDP/91NclVCHnJj1ner/gn/kc/kp3ZnGZobX
Gbch3O49lXSOMq0dmGhT5X+HWAiohS6sNvk/nCN8f47cyqbe4LxjWF46cPII0/JSFyQPq0Zu/hiD
TSGZg2jziDgWa1foa/qyYdX9Qq5nHguJUtqdGko0MYs5sVaXtAxMBsr1WqdpkO8vS2kHtG8PMIrh
dxAhUO/sEqsPtrFJHZ7b5W7AM5aFfcMaQqaODgR+tVWRHPwA+rmSJId4ct35JWQzCxqwA8G2hLx3
yHDUrhq1UjHUILkbXdZusQGgDy8NSBqaTacJiX3rkqNFfMtCiT6FxHH/9Oxp/CPS7F8lfcDRRpyh
KTlC8AsauZb8ejdgxzdXKsCwtIfSE+6U+euAGsjTc1KkiegeZP0vYXSaJEbgyg0XED922xtp5QRM
Ym005IUhsmHAYp95cSKmop94vjvlkU/DeeWRWPZymi9381OlWd47R0CZqG9GjTvude1CAdPCRR5R
RKutlXulXrq4xgWzlY+KcAaUZLjCGvdgj/yPP02WdGLNEPccQvwp49EiUNeW6aTqJldXy0Cnh3II
z6V5P7QkaLTIATQ64POjFEUPlIjlsBQOPtQJshgsi8UpgHKGkH68bCeVf2nFwarx3x+EggkBEtod
5oANMYp3fJ3lNvY7Vu4z9YM4ZI3D5f7ARUnfeuf0Wba3wRZk0J0MmTNydVx0XSqc/lXKQFkf5vzm
a8goFEjcxuMo8iSK+Eux7VIRHrsUhXBP3pV7F46i3foCmGqDVKWrHDHdkxIhw9Oy8P23Foamo6e8
8eDrOwjcd5lE0gKIrLg5w3tKtJPbpIE/c71hnP9zBWspV+ZvOcm5C5aQFi6WYDTVmu0ycCQ/gQoH
z66nS1K5ONDmEqrFVRC/M/GONrIygWNzpL7oslUlq3VkRvbNBGQlmUGAECnYjdCZoaN0j5klYjDg
mpvyKN85wFT6OObm47tFCwRiBugsTriONkRBweBxwe90eWFdJJAOR8XpwsrPWkVBZxUzYQ7K4PdG
YDcEOuIYAgv0yFiEnoIm76iEV12mQ0p1pjWCvGos0Z0xbJLVw6tUZdM5BUHOH1CyjHgNlYKdAvU/
UQcwIcPXndAv0UkYp602Gryp1RiyEKKToiQ/RGOqonJfenmyMcw77ih8x+TGCj2/ySXA3fNLoRdD
XXpF+hQzkrLC7J4H5dKEBiiKxQZIcFPUdHkeAG8Kd2tyg7Y9JtHB00Z94+VcGcdH39V8eZVTTEuW
+a/apQQQ5z5a+n66ajhHVKS2yU2j6BQrkbMDzLuIkBuFXjrJfeTklqmgWsx3CT5ELGKyXj9pVKq0
hFlozZf10kU42DZkjvkUG/dA6bSb2b3R2IDs0XK8Rznfbu7vSbijHLKFYyLCWqRiYFny7KIoD4kq
lCcTpCw4T9woBDm5L7a0RZ0zs/2E8NVCxSzrt+yQPNWJAGQNMqv85GfkYEBLIEwQjRxAt3RJ9HTK
lAQc4mPTqdr6GrtydSdE/5k6dCYahZCbG94nQwtFwSyDGGv8kPCua03etHiORilLfpr6DAo8KHS5
keMZ03q5KxO6Tn4y3iBOM6g1PcleKcyYazgD8s/qEtAHe4WAXhenKtLY9g4LMHgA+QVyP1IEnewt
UuxV97x8cJH0KeDDe3vgXoOQSeGHQgM0Fu+yZ1UswEjesnNpDBNPE48DVZjKn70CnNMdhKg09f8Z
w9lbszYR0830z6xUXVC4FVpxKnhvvKboZxg3JPPJJ9U3mzAasZyoPhaRkhGtdXO24A/XSDvZ2fWP
BV4c3DNL5REZIhVYOcgMJIJAgOLUCqZwDEB5Y8j/ZGHm/2MLHLtaLHQ1mbBiMFLKlCkskbBssMyg
pomSqeTxcOzDvVIFY8zuqRzxel+qT3rUQZAmkceIhiEwv0N3/PsLTvpQ80fDkuVaRLb9aPt6af8W
Mw/nN67BXJ0xRNG3je5pphvRh/wNc/nTMYRm12f3ckIDKeMoWCIIvIvQlQh3jwnHhFxLT5ItQGvY
lGJ7/amWuCk1htzfYDaku8aCANtVPINCdirIsStJ6cGSrSKjQfmdnPDsao76bg6w7LlufbyOrggk
/jBoi8GtQKAl/OV6XQ9tfPHDi9znunW7L2Iu5H8ur9qKXrbh9nwk0Riz0FSIxtbtNFgTZqbX2sYO
lHvx9Eis60q68SUFGSS3nXBqdWjcO2ifjhgZDCd+tzPW3k5cbq1ifvNp5aIQj2cnf6bjVr13rzzN
srgozBgrzVh8OMG4dEE2faaON97cBXid4y9Rj8PWxmiKpFcdXU4ZMC5Wu5UU8AgnZdM8gyBqqVYs
RkdmvoUFemMPZC0QVzt07vp52oeNw/YzeZ1GzA919ih7AKHLxaFLAzYvundPDwJLowxGfNkpNyZS
+nlKKiuko1ZVCo6rQSqRGQlq4ShysJT6/ChmQYmviN+utrNZQMHoS0Xo513l26wU5Zqj2PtLaIQX
Ot21IDWQaQQlX/K//rc8VCX1FBgxi6F7rm/K9yEsS0tjI2Yyr/e10RQf63ddJ4Jf684KGrr5OWBY
9M6lLgOtty6fJqRPeVgo3RuHEmc70U3AQqSv/M0uWdai/T5w4rgeKaue0wHhnTbaeNsJxXXi2FvF
CtH7QYGu1/JHxq4RtSffBvNPbF3vx0eAcHQQ0bS3cH1K3pIXZkkQyqJ8vCXtbf1pzmvmbYLI3ur1
3UnoN1u9Rn5dynHdyXHC+VP/zCzVa6lViQHtGFPU7fWtBOwJ6nI8aHqBXyjHSpGlJSHmNBq/Z4T7
EOoTY6rxIspYdlDe7bC2ScZrffZ9TNrfr+G+rDvH9v6taxbBgL9DLDt6HkEQXZnXZagyshzF9LhE
aMKoGRkZZmnxNS7kf8ewbNuhk/NYTyV5+88+mnTnnTXgCP4JyCTdpBNx5eTzEo3Y4KrEIpYjTPjp
yawN8V47TyhDiVWqkU15Y3fjSvNnMmbaUrcjJiDvpysXcDZn3i1aec9+6moujvq8MjRxobmzDpIM
FauXZJy+1h7H2BE1N7YTOns0hfhNfnKwyEU3PvAzbFCAva63MMFvg3otemHZDA/Vehp58GSbnA0a
pNGtBBAOmtYyiHss5+abnXihSiNtu/MvWS8/X53BTM+WaQ+Sgv1yhcmXEIDbTarqDDbKFTuBeX31
dSSsCPbqt7qXW1rqQ0ndL/Dm8WqEsKOWgZE3iqdPrbLGFmmJJC8RXNhawVjUmtuip5FeRyRC1Em4
h4Jd1VK++emQUvizG2xMsy7HVv7XARq9VvAHKwfA27vWQAr9fAJcQ0zWxLqNqbpC07IrkKw0frMX
i0rI9KSEg86Mq1u+3CsULdvnf94UyjbG5YLrZUUgtHl3lCe6lUqe04bHif2/XZuKZ756dhamV9M2
Fz8/QWLNjaXxLigVHXee7ud2DRin36U7QsJQnrS6zgj0wbv4nzR/YPtaaZMwkOJWUn725hB8meqb
yk9QNlxHHKZ9dbUjgL4I/n0xE62xRR0bYtkAQ7LQpmG9ZpAjiwai6bedb1/XwYSvQQQTEgVqFd3m
Czu3+117m9uy60M0ZmOPSPjZGzBFrnAMOPJv4ngDFJo8vc4KGBeQi1fpghERdekfaut/BxvTpT+g
WiZ6dMIJdap3Bt0nYrsL16381ARXqdruq9Sy9ozT6UBE8BXDYPHsBIGelyaQj0xgdbMsLRyesHqH
ZPvoows/LcZojzZuiK4SPFLZod5Brl5gZhdWD85GMglonzJOKFXnsRdP8d2fc1CsOsREeUGs9+HN
hNnQo3NulCFi23yT0lru4CR+GKqARDmtBQEjbD2vxf3Izy24oQi1dvK6S/2boKdOZpL8X+MJzG6C
mg62FiigljTf53hEBmTMmslaNKW31Qm01+3CdMwHDUHXPoE+b2vjJjcWqIQWZyYcSCmSiMQRMh88
qHfegHWGBNkjNErghsY97PleHUL+fbtIBZHSFN15zL8SU4GgM5jd9R+TQDwk1d/oZv1hIJURSeur
pwE/wakNaJzZojDrp1zBzSpxPkng6k90D0eDZB+f12l/l0FDcT11D91PI2chVAjelqU6W5jAKlUj
4+C7COYTIIjht8Apmtdkk1Rw8OsPDzgnErlog7VMSti72tp8KiFXWR1rjfJ1omVuqLDqTw+gtP62
8hoi9kzTZbASVyxT3JLvaWEn2oJhB+xtSaFYg+LEXRa3vp7GJHtTkOjBmKNrA6Ln8/p0RAqPiTfr
wMipGaUbZAhZ3AztLM2Q+QiQO+xFK10hbbC+i0LWE13qglkxBfqnD6GyFmSfEUP9FjNuH/V5SzhL
Qq6GguNQXbRiiUDmrT69/HuX4upvMiOB0tBUAJNGyEUBHvthwgb6WMvHiuh4nbzjfTH5t5QhPkgy
sh082dNf69h6TOZX7udbfLQqAesLJND921LLhMY4ecHbABYVItAcaVmNmZ+CvkRNBpMmY2GUtHVb
SHv3TPstkvIaR9MVgvpqaLftjoqqkEVVuPLxXDlfBV3hX5a0p5RS+M//dLAGo27/NsxYBJ1i/owa
pafc4W0ETxAGMcSGWFnu1LzbhexJ4mPiWVddv9xo4rvnew7vD5ApJJVJ5LVICfNDDkMNPDYTADQM
35qpwAS8qiSJxrklJe+Nt65fa3jUIueoofpsM3cODGEgwkLGYL/ltkD4q3XreiE1DcMRaUpZNFkJ
vpn2PQsvzp2SE+bbP5h7HHK4XaWekH9ko2M9Av0iejJnzOFRKOISeb7YvTvY254gYmRTL/P79Bjp
F4dQDoKDqVXZ9O/7EW7MYglXsmZQEY7u8uAEYU+UpGOZzDJzf1v9s8Qv4sE+bSAH1aTKUUWH1m2V
UnlEurF3gvX4kWXrCwv+Jq8IozuYzUUYMZxlgFGUWUwG55Ks9LDhN7uwWuev33JoD9iibO1H0/cv
OuZp7OwpQWXWaMxoLSYXpgPk9r9LigA8AXnJoF8vSlI9fwoGBj+RQCHEF9s1rm9625+iUu88ZPkA
V/w2EUa0CEur7mqVWmiGEgXP+tVR2ED6DkZC/EzFRZNSNqqbmDjxEVxmKqWwzOpQbSYvCQNFbNbC
/TWfdfG/1+E2o5yZ1rDyu1Tvaqh1TYeqOFL+TLTTgCx7n6QifLZZwxfkkw60lIjcy7OOuJOAAptY
9vv6/MNCl/1hAWGulTDlAGy0sTvK09kN9ZBWikOAVG9KeRosm8X0Bp3dqBgAqeU58B9hbkzFKplF
2EO/fL8bXlz/V+iTfB+0MpUu+revvPjERT72BbI8dO/GbeW6qSEpZK7JZWWF947vYsdCBghxExlh
TrnESbmxsyJX7yzCskwdLjAxmI1ymNqijqYPNf0OEhViAZ4sM/GW9CEr6NRRJqdZOfC6gGGDi5V6
gNF9g4Hwrj2GdbQOzmKEtebG91/djlucHAgrOdupdgkvGxWukb3km2ZOggUHC/qxFdyhBoIEDMI9
BEqExJk5+aI4rWqw4C6ptfAAhEVQt7In0t3PhEodv4RegY1H5VhpjDPIYYrmbuSOPtlEoeXYhii8
xAd4qZfZrT7HffUlHaYNRTsryrQI9OdXHgmcXIMUCPVlohzdlvi3btqJXVWRXLoxjqo3RIY02x6S
Xpoct+2hj9IRtMCHB8GN4vH95s40Zq78TPbi9G2hUGCjOd6JD4Yf8tp6xiSetZ5je/FRM4we3kJU
5PbzdU4sw/ggC6qI3ADMEv6b7LWVz7J4hogj0YOKxQ9OJgEXSQCz8NDf3jfBr8G05mREZ78n8DB6
UUoNemVNFgyvG6GjNzi0Dk+WrIEV2oYtDkxWkK8s4jp9dRwd1O2h6W57cUJTDUAUiBJ8nXNFthPW
l2/zjcR7VBxi/OYu3I8zO8d4uJ7WfdpU/c1xW/cV7V+1AnHtT1SgXru2zQCZW57G6eTKWLrA0oII
4/+p/07b+Hre5labhtNbuRR3RebptNGmbeZRAP8x2TxVGjTloqbe7ohINFizhA4NEGaJKuT3qc7W
nUE24Uh8kAtAzCRGonFCXlV+5iRcMnVcuwMNBMtX8rDBRtW2dr0hd5PL6nGJmLbJHg+cwcqmEo4q
tI6iPZ88Qm1BCFmcJAmwHLSLreOR8tPSY/VWds8kFJGb8K2Kz4LrMLk0d7L4V6jcAsi97xnTFJNq
YPOZ2dwahQmlnXAz1zNS5IOZPYoZgjTXrr4OBkAVMC0K2lb32VbeLQduM+8I8d0y69Wz3wBHm6LM
OMzQy18RLnc8HMo4MsotF1dtaA9ufu/EOeRwtZWfLTZ+nFjkYCCn/dVlEIdf/Gd7BMmbixA9+mJ+
VjDgDGEnEEoLmYpGyc1BRVWGTMALLcrI1EbCq5CkELC1uRIpndX3NfN+LfMIUevTlgyCT2OIsIlC
KZ3b7tMBn8mmbCzcoCyHI2A8/K+YGfMyf68DeZY2nkBm3M2EfpGIAcqloF7nfWedTd2FpG5/DiF0
8Q9WD5oWt6Ii0fYoHQR66SKve9uR1jDYD6gk1jtTNN0BoZHmziY3p+GWLmx0QNdETmBFB+OHBtH5
4RzB5kIiBLy+R7KC/Kaz55y3K9y5Ulg+mh9JAVRbJeAJzeEGYmSarfb2ZW55myxmrWWTpfpvsRR3
Rl6aN4WfKEERalxKORkeUn3alRjGelZq2EEuOfD9eejuVswevfOnVFoDQlM8LNjCiNiyFXR+UgqG
fe+xtLEmCSdgHi0ro9yk48eaNg0eX8j6/kWYYKjP5xf6uj3FeSt1aDikFtxaprYLxtQkRLwAuy5v
IzH5typXwKeOq6utnL4JoWaEw3qo4q9WJR34Vq6Ehg/ObQ951Z9ERZ2VB3lPMt7mDoD+pcmxenDK
LAJH+R6rDKShGP4pKlpVu42Yn3zWDegxtl2+NwpJrQJ7ZO9gmVHsDhq8qd7qgox+U8MJGVnl+P5m
BUNsRBB+xyCQ8vek5biZRGP6p2PMCoauiOSCixpvXtgOhQUBl6RuaXQ+SRBwSRhQqT3g3pQr6p4K
IKr14gavN0OpXiGLGuVPUwIpqzmXLz6ghGVMsg9B7Zdb7+w5T3UgcbzAmRXHxEbMpOy+upfCRVIB
k42XR5XjZ2UDs+8LiplfIYZ1V/SfyVqhQRX4fafViIb7kQMjWhAoY+n/3Dwa48/iEjxbD23lFZPp
kYUhilXWkR1dOJ69/tOMPAo2rwlUYfH+SniKdBuBlVsWIqd4xuQCpwzW7SJkClE8ZixiWrj9F1ft
9RFnrJFZYepS15owajkLZvw2fdpOBFo11e6IdMORHDmLA41+FNDkbhYLSh1CPOvF4jpyUEKuEl73
kw4ueVP0h6RnqjB2UjiN5qXX0Rvk9ajgYXMXYSbD5BbNSoR+UoB8fAFoixfQrAFCYCvG6eBdP1GP
5xLMxPdY42YjPJvnmlp4RkFKAp1Mq6uFjez4BA64v1i/QAO9JZA9jNvOPZbN3N+AvgmTN1yzr+/z
ss6IT+gV68yh8P0NO6dmtDtcajtjJ5aq5oX3dS+H+CJBsZMzqnTuQ6z5TBqZAz0YfCUD15yfEc4t
y3xhXZDC5hOc4sS+uRdnpOoEIJUNn/Hq7fw+k5AtD3eed8AjUNWwieFVcVcjMxWY0ksc7IfK/6iU
qnu5Tt3KLmJEymxuTrUdiGHNS5p5VAawkZYTNANMCY5BLMQyE7uP2D65vk1QIsU3B4QD552j7MSn
bZtx40NjrsaHZrvhm28f0+HNZP0YoYCKroc/X2OP6m0IcYLa1QIphvf3OKONPdis8MVk66jqjbAH
B19hrGHorx38QOzewLNKCPoDcVCgak7UwtW8xahSMF6wRWOE0DY6PtzXwalKv+HOUbPHSNZxYGKf
ye92zFW8izQjv+ry4ewLeJIGoMhlNqC1aVIuwhPalD93UsBjV0bNEqMSaCbRbPWpG2ESapdjr4BL
WPSbmVGO9ps217QoBv+Mx60m7sPjxmXFNxdYssS42NOvP+wHMmG5B7B7G9OQGlE729ZoVLpiy8Df
0jatEA3eDBn4TyT0hzkmFVX0R0WrLEHSdE/k7JlTuPalBbr4kXO5VXc00TqG9fduN7AQSMlmm6x7
6+O+u/gg1KO5euvgiwGpEa1EiY/upqHcXiM7Z0VlMZrS9AMQOquXWPhUhkN9fQKZsiC9fz7DA+r8
y8r09d6QbDJt7KKpcBP9JDJCqA1//uLsnEJGQYtVJbcyKjaJ7bL4pEMLma/LfeF4kRouDRVRSyQW
bfyX1PuDDyrvDKqWd3djGAqNoYVGiPwFfnyW+g/I9Vd0zPh/359DvLoUXxrSFSB5Gp/DxrEHWDeE
ukqbDDToiANvCOKDZ0uyZcOS69ZXAE7zqIc0ahVnofPVYZm2SFOfR38vocwwExs66xrrQMFCQ370
LLr8ivbmKfZEg6g/k1Vj/8txh8uyN1saxlenIJ8s0E1x2o0NM5YPpRoZMyPKWfdqY/N9OW1k7vPr
7NnOGKcJ5aBVVsgrWHv4OTLdYYOWgEz6lsQQkxufCSEFNWLIbgdpGXIP/5DJ/BToslvgejtalba+
aPnBQ1oezFlresxV+zp2vU7C9OMEAb34stRLE1z1/utDth2Z7WlDMBnu+9Ey8SluUuOiZiKhn437
04HVxme56ijxIDVNZK6UAzHNX/rmi/oCvvPtg+5+PjLdC7MrYZvLiZ8rXlskWWoBWl2BjfB/KOdm
PkISWEWnThyUy3ewtH7Nm5LFs88ljwWcKFLfQ7qxk/klXnply04kWWSF8O4Ga5CoabPtXrJxp/U8
av3KR9L0JC56/w4iY9wSMO3EEMYIpNGfRipvzHUcsbPkzUeVfcRUiE8/ihvvJPy1eWn5bCB8CQ+O
T1lSj+FbbSFz5hHLC8SQxdHV1SQgZ0SJrsItsL8X/pYSYdeDS+EyRCNdrbdI+lUV4qaBT4dPnYok
lq1IsvlMgemeQv8Pb2EpdKf2Noys4rpT74qBZlWm3BDbY+vouX5RJCuhULu5/LxsLYFn2cihV84f
H/3CWJzFoj5EAm9IEh7V1dHNRjTo4XV6F7OKSOrXE7Qbeq9IyH4weh/GcYlOKj/EGbtjMFuTmsmZ
FkgPvr9GjZmr/BGAMzpz8nE+deLDYsmfdhDP39jHLNe9XnqgSQtp+/NuEsSU8LLvae6r3Jlx1iQw
w+SDraCMqKa/WmOq6OS8nctRnjhfMszQpWir0n2tg+Lx10q+sckzn7UrJn/tFzTY7LWQFCGCdxtB
K6RihtTaNbB8nH+gFHgOR8+x0kgWfEoETkOJpPy7eod+jVuji96k1wfOjNAXKtq83+HZBqlRiBko
sYa+GpinGLl6lxMHsLuDGA1gaDffbI6nIoYEJSHE5cmqXySGY5bAQfAohVb8i+lzg2ChVJjMiEmo
xPNduOi/euKaj9bzm56T1zM14VbeoEANhPuMMCf8Kq473H8VAocu8Hl8rdFhJAkaN/ozx5VP0Jb1
3tqf17S6xDORl9e2jR1TAY49eMvHEdtdyFojp5ab6D3LORmWacXLXUNXWng6r3wcp1f6l72BNVZB
uNQPXed9b1f/SalFJQZuShFpx4H0t9Nm18+WxHN7hbZCURqyHII6u5jN181x7gq9OSjhc6uiDCMR
VzK4aZO5nE0+nJESjvsnIqtlDgbARkcfuJAUE0S6HLGcpOrv6jIHO2yXJkqL9bK4TfW+kAqGD3nT
Dwems+hBg5RozbOLePl+5dc1wKUsW0NA2/QPf5r7UrN1fwq2cSzfE9XrCdKf8723qlpIxqmSSfs9
E6CKfzyoEM2ANr2qd+0+hkyzewdoh9MyUwUn4j8liEm66eK7vrf3He5yhpPvzcoyLE2PkewfC1QK
Rztub3WHVwHwY7VC1JIUqk16CqSCccJJ3szOVIhzJa7e3ogv6bwt2T1NfVnmTonCqwSDu/mxzesW
QTsQ3zWX/y/0MckVFoK/PK1xw1V5Tza1GQqpVLefUUZOw2e3FZGtJp/9p3ye3h7LHn15wH5ZdDWK
5ap89D+Nwgb4KLdoGnU5t0plytGQ8VlZ0JqyHmzwV12Gi0HrSsJaY28+jn8uSFyLLVbVgLjvI3zP
WG+fhe1aatt92HGkOUk3b/1qmIyHe4Y553JgOAEUY82H/jThKeiH/aGDdju9GLqTAJkevIYcO9XD
cVr3skyoO360IG4krApbVtjgQk7TM9fQ2mJuyR7sPr5Vrfy2Ix+ckllqjgQg0LB8ecAokVJUQzac
lubMugKU7/Ix3FxKhQHNwki6tgJxFFzdou1nCJhrMwSz6fKfwGccY1OHY9+whH6bpg4MYJNXDTqR
4N/t+phSNkuWCzrLuhHhcAsAv3LpfhlxoPqI7W0+DMka7pSzpGpziPC7OmGZu8bN0nNS9XhLCIZd
MVH72aOoLTPtxSLc3DKjvtwvRUuH3oSLlppOw/sTW/05BPniKQZQJfNTA7fiUPtQw5XnfQx7BOV9
OV4/GswQzR/o8PnzrDyGNsBaQRnLSGBX2rT0wJQZogLm+k4/u4z8igwboFk6M9c96OvwaAQG5SL2
L3XipMzazt74xPYiBkxbdDKaVf4k/aJ3tFo8xSxqDPviFBi9Pgr4v2zOgNAwgv6s4CSTpiogFPNS
O0HyutM4MF7qchrEBSncmkV/Ge+Vc15U5EHqoaVJCUH5UMLnVIKOv+ZK+Ga4jLr/ClNX5J82xfNz
WIEOa6X5el8YfYK21uL0lUuHnJMrqzIKQm/q5BiWvfEjqkWBCO+WHXf26+mDlk0Xx24rVLJndmcf
zd5VN276kQ0F4yJ/hgDOwlUyDY1/aqMjn+MinIHBsLg4h0QOpE+cV0HkymUI9hVdA4k/QiULUP1R
xXCpU2Q3gcDDkdIwBI5b1v2j5VH6cWkMt/KUDeboz77QwEHgstqLiYXTuiuA33zKV4WQUA/5J0QV
g3yihTBvhyEzFgoyxGuK81YRCBxsAwQ7z/d0tWc/cBRGMlMuAPdpFepSTFXFbkCmcIqmIrCrJFJE
NQc+yRBUCxzYo2CPHRIJP09xlX42DdT9ryaUAneP0s1r84/TPLaFsMDmWfo5BM1zNGlwxLZZqxiW
pJ1WsPYx3nh1DpZhZVdl4AddZW66WdGpRkAi307Xor4NArgShw7kIjN3HoTXWH+zs1hSsJf0evxA
K74a0zrLzFSnGy6OA1k3QGiGRbSOJ92IJdDk6dO2lLWrCapQkzgdtF0L01YQRal1Umfxepmkf1r/
czhszSkjLdLFq/Ikk1ehC+N9DmhU1FFyimdoQqMQ/zRAER4KuvxmGXVfM+ZkQMPVt9F2UFYCmb5n
GCgzcvASVvS+MIDYhBK/x7lJRDW/APY7X0C+JXz/KoVhQzaPOrC1VYff4YhvGQLKO2GxPfHTrtHI
sAtze5pWCjcKtarH2XM+s6GmzA5zMuGu6wtN8ycpQ5pQo3ynbqzTgPAFkTektqrX1dOigVFSae3L
SeJoUpRatslD6zGg1VAnviLEqpwWF7SrrcNvYDixSVISOAdncYC35Eew3Jfr9ndAc7pM44EjchHx
MVPlDeInN/6o6v5jMONh/R4+6Lr6Q78gEsqol7gt5tcjpnwn3AvxzZyJ6XL9ULvQrEs35eoRvkMf
tFbLv/3a0pmlBXJPHtoOxCxr3JhEOOiItS3XcYlNjNCB+CerdCyZoeU9Q5tw9GAM+0m5jucnKa9B
QaVKCziE6mCzVLOf+t2KWLtyjTKcxSHwNdTXiNuUXb1QtRueNDnj3NAqaZrxDfi7kUANlIFlnaqE
RGmnVyIu5NJhVMWo+SJUY4SbxSzPa3CA1r0136FAUZ6XWEgFlCANGi4HQl3WoR9W6FN6iTZhSDhN
AjJsZH59yUwH2ZsKvEDS7njtLbsHeTj1O0PUv3Im/87YlPh5T8U6aEBPX4nafYmQBAHPaXswKkyu
49cah30S9B2dotwQGhyzz0HbQty4hrZoPv9SPFqwao8Z3ibhQl/ZFP4FO9yxqUSRigE5/ZztN8Xk
3K8ZMi14HkM3a25JJPFzM/CozES1jlYgb08JOgkb3325Bp8aZoTg/1wQsrK9cKXSWhbgklsVQJP+
B/YDue7ebZ+uuFfMeqzTjzKA6Omqgq1wOJtg20anhEZFDpB7m+Dl+8T05/GdGj5SUkvvBQT203Jj
N0tykGNQqIpQxfFRRwEL7jiBzHIxDPxPqP8aF7iEsIVJgBsIgN5GYZPMZ2VlJHui5aUwtG8pu7yf
cA51Yg/caOaRnW08ybnxyYhJCH8aXzHZGafaV0mqZPz2q5rpyN1EX101RXRz4/1TV9GkOOIfzDaZ
8eoxVrMo2JO0dDxn8NAgIDe8+rGdRVNzS0WqcTMpwwxEm6wR+BFZT7n/ODJflHlrfJb0Kdk3DXXv
oTrCHbZiGr5LHbfKU5uYXZdrp96YJn2CrqKXGbU00L8I82Q0Dm8x1IsG0GKl/k6KpcIenrCMwMVg
27FHRr4d8qvZ0sduTno/4Q5aCvKbkq6Q17Onp0GOM2mnfnMD79ZmlUn16M7QcU5+4c2DcHhK/7ue
306/FnQHsVaxFBn4vFalD+BIV10Kc7W3VN3yadZUKjvKHCF91ICZik0fooOofuaJLzZsBAZpy2Xs
v7t9SU8jEBbnGTGgD1TTZitEeZ04vCTtPn3G53t/3VjEWU0NQOViGEDNhhz2kgVaw/DvP3EnYftf
Rr1NNvwrjI7A0Pifmi+4afAFwrtbx5DkcUdzsrkYvo5aqA/kRGiPwfT3sHosddrQnS0WjXLzTQx0
GtKXlOCFWofbfO/saWknjt6wIxcSbjAZPxHi6J96TwCbRRyzUQ3Jc29AMW8ipjcnOdGhMSzkwWCd
Z42zR9q1q2qdzdnMGGIraPm0+QSKZQwUjB8Scm8jp6n54r2YK0rAQEuGGp+EECJnbYnj08tWiQvQ
05g7PHPsnnHW1bQsFM+g6Mp5HtHaQn0wAYffkZGDQSrB+AeopNM7UgZZ6RSGBy86iJ9E7mztLxS0
FSkMWAN9G5fO6okZKfa08u/6vhnivG7u+O/ei1fLjQWi5mLtStReP0OlTfs0uC1qNuS8xVC9PtTO
AgkY5ezFOiQH0vwrQlB6DVpKbzY6O2zHgwDgGprGFa+p8qMh9a6dCDlrr+0H5x/d13mpYcdQkFST
6amavxQQCPRqag/FfLITdhZOYrOWY7vd3PX75HWk81r1TISzPm5f4svdHrbxwPUFeZ8GV45WWv8n
LXxObTSTBBlUdJOq/vSjxmqjjPjdpmIVF7gkEV6gWhTMxr79no6ODhvSChAraJNxtx51kq+LPwd0
eZlT8mThPjMcEFQvfY9fsSJNSxHX2/+ZH67cKraVxpgusgHXdYs+W8pD31XSN3MdmYzmDNTrDgbh
nhaqlaCAVR4N0iJq+1wlgPh1VzDb+8L74EnTyQvRhGmPqfPWkQCk0cKVpq7gjtJKXudNir2dyQqt
8aqlkNprSNfZk6K/MYsfYiSllBbBbl/UE9gO4rR0aR2dD3RuG4PlVwX/oy9tHZ82n9DWp5ZsRAnQ
KYfb2w+GcUY6xxQjdrNZ85P64/IKu/sk18WI0DG1MXjxGtjiBE5F8oaBv97hBINc4dok28LGJ43L
UPLBsXfNHHCDujccoWK09a6WgczPlvOuaCNPsGlkzedceW+nGgD+pyDi6j5gSnw1o2oKKZ9/GKd6
9rfKmIpAZvN0sq0VWU5RV+QGoZihCNjwad2X6wKjayspCxpEX6FtivQ4+KIpcVqwVMp10XNeXbC0
CpWVWmZtBDMeLLTY2kUEJOtHapLXhz5ZCugRaYmA2d15tYX69GOgYKN4zvjF91d5K8F9Xq3+hv72
GiEchU4ALQ8cJBzbNWZ3THJ2cDIL5sgMBU4qckd0PDXp96JY/kvvIqhD8ifCbjZRKAwFAmr3FhwG
KUreh2GyJkjDvusQ6LS+5Wrs3js3jlGwIrU3x/lR7Gf7u3a2lWQKw5f80hulJ4X9br1Xm0yS7Ljm
2BP1LFmVPzVF3yqMZYajeypv46gqFfwlu/Rksh7WRa9TvCLFOq+C3qBa52KIAH7Wee+v6JZzdBeN
koG+W1mZxssEm2ibsmNwnoXS+JPn9EpHI6E7+Y70huV9iSkpupQJs7VRZLX/wr29D5RPs5/ia6DN
gIF3NZaqhlbruDxvc3rjmGn7MXJHJO0cA/wcBuZSGUmAopJrwIzMVtqDZkRl9qMJrXZLwefLnhup
6tDkf5EhPa70y2vsjVG+Xg4errw2fYTuCA2aiaVQmPcq/Pn0kD1O1xMI1/y5NE7b5w9Y18tvlm2k
vCmtzRsDFIXuBxaWDRl8mdF8NJx4CuEEOcG7JtPq6RIceJKa92rTyAie+alDde+OyAYjgSsQPQ3E
hWbsWQvVNohc+f37zkmdoSPvoN3w12+E4C2b5VlyxOsCLedlTQqYUZmvaPKSdVUowJUsP/p/Cenf
96u4LnSkZrsmBvqRLgzAwfkHUrjj08C/NWnovC2rvy6xUHanMyJ7xTQbPzVmx5fGRvqTkP1sU0hm
EOWmu9Hnvx5zv65QaL3D8sw/7yQSUxoRD1255R8bmqb1L1aAoXKWJHmSGiZhjIgYuUXHjG4uyBw/
YaUHTjLTCjm5ceok4gb8P/dqaAdNuMFFJ1MTRpOqYE8/bJ7p5ABTwe35lAvtcf73p4QLjVhv2sgo
bpvUOlCic7RakjJSvXvo0XnRzcpGwFzkPqiDH5w8NhRZJcI22ARDkI9KwqkBgCdCNqcSTuK3IQcw
OwgUZ1+/PDmEx3mJCbe/eI+51WXN4hszOBWm1f0aJ1pHPbQQX62zRsm/ZDo47a8Ge7JW/7LQZO6f
o4uzvOOrcHJdWCxdw+LGWs2Ep0R0at6hAOFvSouLZVKz5RV1klAD+e8i7NyKDKY++PX7ONkLuVx2
zUGvcwZw8i5JKfIvqE//URH0X6u+GvrUIasaWDc99OVHaJN4P8K1UcesplxRDp+DAbBjdlBkzNq6
QjB9a6ycqAo3tD1Q1l8U+CpUcO1SpZdFQW92MuVmdqkL7AEVABhIb6SZVSPgeS/BoMilyu/M0lnU
yPOnhc50dGVWmTaBayGtO5sIWTDiEvo/gfSlK0uNc9OXomrdlgr4EHcAUku+OhOTQI2mtepnvmQW
9zHMPyDizA1UlBz3+48PiU0xDva0PakPPqrYFZD+3QMABKsd8CifV7ItS0/ls3BfRP9CQ1i7Aat/
hA8y0f7U3xLBYHDzjuN7mfA0r1HLmOAP179Knse8XJUeB1AhDI0AVNEnBxhZ3nWFYFcob6wppmyw
DnBIa7on4wPeLdEA4TADXDBFXzur0Or8SCwynf47OSWcLJyQly29wJ6EyL7nZ24/C3zdUYsAyvsx
dam2xXRURk7YddSG1d73Q7fB4Xkxkiele/7F+MsFl9Aau3RJrqe9CDjr1ALOl9J2/hm3YETeTY27
w3ffsL8mU3IRzuvIxzzHX7V4y1MBPDxGFubC1Y4mN8ZtMZg/GFnJEBS8rTKlgsRwgwzRl7w/NEoo
fdNWyzbsa0K7yQ6D8YhDHwUCWAaxbe/0hjpmnKIC+zEZCtTrXofC5EfsYqxQQIumecxC3IUZ9A7q
oSl62R6mc6tnkB8Z+8dLHDbkfPvpU25v9w6CsVthKH6udCy/pohH23kcWJFeAXdUAYdK60Z6bwiZ
Jjqh/omeujdC2amIkstPkKvUdj8YsdKHywwsLPtE9GkCgFGWNOQ8Qhocm3veqwm672+ZYU3viDwA
QFA/QyCEm7cQiCeJ9A75jdbs6h0To70zrlqcWB1dDrTx7ZN8ljpA5T4BhwAHb5QwUOs8uOEc+nF9
qoPB07k9FLANP63r2TeBD1t2LDomjLK2aCxplXBuBYZ5doyuqQB/6XzIwC/U5H8i629mvC4m47Mj
PaaDN4qS/VGTgcQFKKckE8olx2z21+7m0Mblmp3idQHSkY5K1k1mQ5qPRsiGl8V4sjUwlXiZoKRK
yiYAwvSdXTSrwgo+6M3uvUMafYML8yYBw2HKNwxMrYKYoFWEYUSj1L+zKMgEIePxpIlnC3eoTkCx
0LzdkC7pkeuSb+J444qWsugt5uRpLktmcJg+I4nWWxEdpANcfYrEmLau0NiZmidY61/Af57VK9aU
QxgEH09o1z+0CGhOVSM+pKcrNfHZlMa9OE5ZJUuU0MvRTL1Y66MkA7Ds/TRbuaetj7eChkpMTqbh
BS4/LD9Vr/uamfQetjYPWUGzlELVCW2GAxpdvEDFIAGIjC4Ry8XwtnLq6PiqIMe7pxBijGcKArJO
Q6o8jgyZKUv471xHkK323EoNEkMZweBUApJaDXsUafxKop2Yw6bsY0hVUsUPsyxkH6GxohBi2qp6
6Dj2c7+2xQE4g/XwT8fqoXvHjRwwRbtYPzRFxVsZTni1x2gF+4F4KoDEXCTFR1LzAZj7ftlhF/cx
ZhaDbSztpctKErn0ZW7S2RvLX4F7iaQfVsBAaSl2RmefQWCAzaVgxfrsqIE+mEJy8uMP/zhb6DGO
6AcRgxRfu/W3ugzGo550M9rBnGohj2s8UyWTzjFU8KcAg4sJQQ3kinq1aar9fyxOT3N2O49FlusS
OgudqVRGfqgthDzKFqneUSY3T92vJ9dyQ7C94ZYxLh2irwHBPtS9bEzyanbTI4/uvy6Q5UDUVaWW
7k+BcDiwRbJnD+QyHmBPfhWyv/ajhrit00neAbKxmdTjrV0rzZOnNsGT/dt3naIAxn59poqnUmpm
3Ukd6y5eBDh5KN8gReDpvd3Yb6q3qWa7qLXKKGh8OytVxa2Se1po6at52f7bXMy3Ezwkff9d9hft
ktfyzrrDGb9seLtH6NOlvFezvJZPHOEs3QKNNbwFQtgkUU7/PPS6m7VGw4embP2e2uZJJ/H5v8Oj
8xRPABK5htcAglFIENAG71n8rQQANxIApWpsiUCx77H8isW9GF/Hk5ZcFqAFfwle0K42z4pwFHW5
R3nD8AQPlQeVY5d07hdpnRWDc7cSRVCAVd+hnXiz5kim+eClq6CmmoZsKoW2+x6hEv6ShXb+CNTC
nPRaJG3elZP6dxvUMBHxfxTd9q+JovzkAuQQ7pL4UubpflSs33XwmwI6ceQBojQqYdO184JprEx9
rl9WYKpo0VrLi848048MCKmiLdx3NlI2iDUdIdaGSYn31PDHip/aqETV2sg1JUfihnpB510Lgdf9
MKhJtHG05RNcthWiksOAqaw/T6BxR+pcYm5+tT7DCqatlqcHV4CIcVPYHVmB4KWh/7UfFTkvUgmK
5NlNh1W4tgzN41ia6PnnVkCOKpoYLwap0l6uktv05JZkW821kmGkQV2Q37v+6qx0HcqBUFl4iWpP
YgGhaAwjDJ488CdztTSVbF/ebj6JkrG48XgXEFUL6yM4lRw0ydA0E5xaZgC0RNXfeIM09PnISjG0
tB7Ed4aOu0gCxycgq4N4XNi3g2Cwjk7fA7yp+MrXNVHb4kEasJ7Rz0u4ZyxkUhQrwvcX0X8ZpvAy
WRfGd0Dstih9qF3f9rnforrZOyyVCqvYLYBJ4nFonnb8CMHuA1dEpW+JFOxaL0ZEewoUpVFGk6HX
jOL9KtKA2aMlIhvQC24FAN3BLONqSZ1jGcRsO7+I6KO96pFv6Rls+Uhf1u5WbLnUR71wEHHL9ALo
GouqrSSJazbMWHd2ql0m13vvfihn0hdNwDQu3ugvVElZVH04f4Iu0JJALiqrEaRc6q/jFXM3f7RP
Tuj/DDoPzwrOfNEXEzY46pq4Ft+J5cY3U3/CVcHJVeEcNdSdlwFxImAquBkD7W5D2bBsLSKFSNAA
RZXcl9MuXIqkf/T31JJj/llKfT1LjWFeGDpk+cth2p0Po7X6j5sDL9jIhgs4v8ZQ/TxV1PIY425y
v7QcKKYOILmrFj9/X3xM5cVFQtOZsVrwp+zIwn4yIIgVANaRElbIoUHENFq9BU5H4oKXVm42Y8MA
5f7uIXP5AdRKwajSGfjDhfDjk9yZGJ4qxY1KUyR5PLRGwJhmOSy0mvtQSEDPXhOFTyj/NqFS3LCn
KSXI9PjujJb6EJrdE1Ev1YpHbbM6aF7h/iXUCILOjkgDskSOTg0JK5ivgMy2opHChZVe1QSoFWD6
GAmeiM85f6yJ7O9Q2kDXsW2nY/lOrAx1RCTWR+LQI57g/EIrU+6fFnzHQKs4dCKpkkWYF27b5aWi
XsNSZ4iRzdBqaO85j9fJ+NgumjuYfKZrlY8vZKhwMnZhXhjig1Tw2mJ4548XL8rmf76OCRIq0nSL
hCs71xE5kAyhDLYTUGdap6WD+QyuNcZIrlVIc0DrhEgdIieYQu6CMVLK7ClLcNpeSGfKQFrN8uOh
AaBD2N01spQsc9vgK9d1OiTQTrSH9Upfqy/9AUNf7OttAxAdxjwTDf3Z22qOp/i0Wai9EZP+1pgE
DSmD6lwL9zWF1ftqguj7x2K41BOPAzpXRIdTRlRKtOAsq7g6sTMr8jofPNfn4XKmLkBf82etp2wA
Rmrie8HSOMWi3/yRa+HA0Of9AnxVJazMt022IYPKdjUavrRK3kYSDrTmaAafBr9wPrzQBLRIroas
KOKv3FO5hVPN4wwAO60+xXsiB7t1SQXIDN0/pYtfVNmHcG81DfKl9X8P4zLfMjYOJHf0HYRYw698
rP0go0tGR3+YBiCx7mGn+PpxbevAY313cqdmxVRhLlL0vXRd5oU2i7LTR/VmZUa8Q+cxTudWGD+y
EgSyuQRLZuFQ5lgV7OXQoB+Ble3O1YXyEIQPcjwmYN+ZjP3MnNWvpNKqgfw5VMpokAI8VaFXzpm1
dJfFwsNV9pZw76a8hKOhEsrnyoC8anarb3TkCzxWYIcVzDmRHt2kIRwF7202ouaimGDpeGyuM8tr
zqdzEw5gV4Lt0Z9dOygaAzdGkS9zkGkcGF9cOVfj06i1J6Z/ny5m61I83Nrx1wx2evHDTT5CU/dt
vD/1qRl14ODfqlS70YaOUwZgP+Wj+DQTPMn8L5wd7VWKYHZBARnK31VoBuL8xZMh0fCeQTyR6bGX
HIuNjaMTe74eewDE6pBBIxHkhfohtJbPOpQtENo+SJPxsVKSC/w2W8Uwi11puFPjwMTMf8rbS3Pt
uJsvSKchuWi8inb1yZ6z8y7jxK7F7yAJptikamdihLcf8JASPzLrKF9of6OGLp/1QEGY4WDUK3t5
WMl1uwZc6VTrIkWegJv1i5MuVVmvvRLzavQSl3SBm/7ZnkGIys8hz1/E+NcUq3ObBmhpe+5k9SUz
hFhzJba/g0LWYkcUW+hnU/0Y3esrhCh+kXLliNpTIBioXyG6lr19arOICd9beYr9i0ywPGTGLCbw
Yc25ePlL9CuGy0m51Mjz3DAOHgEe0m0Yd9F8bEUz+AFoW1YhPBtcBIhif37CVM0s70mYzSb3IjvX
PBbjRe65hXYzzNF4f1PP7s7auj1LovzgjMqa3ykPdvEuGoEXd2Pyhc4Z8jiTb4iY98p6HoAGK2Yj
Cl+iGauiRT+njq36svQ+SaUF2rha0o8Q9f1LFUilErMT2f7Wr1rlqkGy4plZ9KoMQ01Z2yKzhHEs
hfdPuGbeEDkmeiqqYhfl5tdjP6l6Tngy8SXhVHWxVi29Zploo1zOQ8kJWShBmt0jaJ6blq2wQe16
W+M3e06QJsToTg3em0jNf3CLzeDUOCiPccFObDZmzKtHpiLWDrFrJHSJWp3YbnYy0R6S9W6ykv6x
xPwBREaWrrJy+vuI1p9M6Kkl/nxecRkq+2Wy432HKbUhla+R11QeDSUs4wEDIuBLS+wiwC8nC0ir
yuYs3q/hpKUHzqeGWn7Ac98IIfy4uzu9FmRprTghpJtINsktNaeFul7ZAdyz8S44EZIGkSD2nth/
C/Sf1AR05ihs4QSVMC/Hx1yxFhYyFrWHpz7LTfNB6UEV2ZTWg+PEVbidlvYheHLzf3EZaeBCoiTM
f3ttpAAfVzKErhMWTh+nxEdGU0eJVsWYNuUzmhk7mtFvF/3qZR7JVtobZ295Y1pJIpDelVnDtxmV
ZyFH8Ekd3PAQpH19z0CtLCQFASdq3/73FjTPY45daeBh1/3r6+RsMuFpxjvZt2p6z8JeLSAgueMm
rhR1J3JWf2Zl8PxWdwZQchFoUne2B2rr5KObs9Ozlhq+MVR3XwrdCcrucRTCukHEFoAZHwaLA/+E
rHdx0QWBAaVz9h9sMZu8h6SieseC0SVCoMaLW0TxssxbUXm8LTc5IavK1oKchcSKtUrycRZ1JAIt
wnEYLI+1lbJPUGvLYH++cRjY6WFvXcQe/+KYVy7C9XGrRsTVDBOBBq0BEN8epx5Wp5ZuzHPG00Zg
zCRP/i89QgMvdGk/jSluqgLRRmf/Tq18IAYej51QWJmUBm+e/q//F6Dj8C37opLmH70TpbLIGBw2
diJMlPNmSjwx8zxUVO6IVYv0oFKTp9JdnDjQO7DelRKSeDn5W0Gv8bxV1vqDY3itnoGvlE6QrpY5
PwPvLY/Rw3nBXiMebK7pjtgbQ+4k6V9SPy5Gm9fduvXeuAY0hij4X4eNgBaBM0DU0ewB3UlbqcRi
eXzFAcxw6TPad9r6HXLI25Uw8lzqELW7HIlFrpFgKP/7O5jeJxinfG+z34/P1svBNIWXzOdS8GhM
7kG9WftvbhZn8IHzRlLmPwA6rjNpG3cw69WF9IGx7KeDsAjBrk977kAKWZcYnf6C2NyLXnGWxd5A
yekdlazD7cAqr/8w/4N8n1mg31Vt+Ux9XT+AX6lqZExat8381ZEcF0Nwn6uTi4BuKpubwBwNvEKW
B/xaN8BpoMqVAgFJhM6/t0kkX1+3xjcH3gchjKW8XoooQOk5E6nNaYLWMLB/UDs9A2uoo422hAzm
+8bvRv9KJgDmN7q724daFg8FqitLKf8dvQe2fXwBGf29FldOk6mqlNve3VqG0qiUooRZ77yVf0An
pDMH07REet71z2GuyT3L02NB6cr8v3V1z/FoglovPyjrfVCJp8fswdrclqvl6BvneEMdMnMVkCCG
EDm4XnIjmr/WYO3f7fDn8t+b2K0oVmA/BGd9egWp0iPJpdPUGW2241/eEqPeKweoGoCIzUYbR0WM
XP2GE+LqHA9KSsW6NJosdk1GsuNwY8BnA0kfSz9NyqiWolimgwH48w2TeeyAffyntbWDf3/QHJGC
CYYwC4XnJviU3jArdHPS7Qw0vIXjTvymyQOOshc5BFOwjej9inxPcEqGamGQ1KEHxpM7W3NX0JT/
MtCCvOBkYkIMqrtt9mTLFH8Tkify+dFTD9Z9f/IIYSTxwjcHoCk4hkTx3VEd+YUgZqOWXqlg5IIs
Gb6C+4v0nW+q7YQ2VqjqGZN33FWPCrw3BNB1m+JNoVNoHh4KphUvXuyCDrfSL+mHPzVFBLHe8oF1
sImFH93b8eqGs5kFNu8f/xBXL3aNJ6olvjIhueqTzPze6Gy9bHQw0i9SK/Or76rHo2Pq+8pJkQrP
CHHyepBgT44TDiA7aJa3Xp2n/SbS/pT3mAHFxGM++YKqrpPx2STc03PnE4L5ps8xdhrGEjDGYQ8X
TYJJNjgpXbUTmtq6i63gpvqE0dNtQ4qlnin/I/7zfu4L6RrpUiMg0pR2xhiT6UD0YfhZMUR+AHG4
DHrCrCMAvdG82RtBZQNuohJJyoDMyAnTdtu6eQHXDcMuyV6IGhKEyoug1RF/maCL+TVuDSQ1W8Xw
Uf164gdD6XofsC3iNHLPy8uU4oRd9Oh4Yj38vIJXZK0Q3D2Wvb9v2BWftN9bbz3ht4B0OIpDxOla
S4Vq/dRvQmK4SpX/m4Pk7mSwgewhWUld1NGautAx17JCbBYoIJ71uWaY1e6w6BW5A34/cmtx92Q6
bJxSX6sT5LIfQO2W6+1wbmWDmS8guvR5dgMVn8FushtNl9/7wurF41BVZJ1ON/xmmr+rdckEMr4s
EH+bEM3kduBxu6cgH08vQhbaDRZjPDb1LZgBeIShxSMqJgg9ioexOpowbVitQyw9pLZ5ugWsBLge
q2Vvk38ozYvv3pbLi9S2gDMQQ7vmD/12Wdz4DHfj3f1/jcGjRknVELxmfQfNzL2W/SEl8hGbmH91
7vIgVkaMGpkf0tvBSi0L51u63UI80JUHIiq2cHrhCqmYjajnJtBR+45cjfO4ZK8ybDTQdpIrq5RW
fQDORurFxip0RPcFih9X9Ek7WHawAjlV8MUkmOFSNdCgBQ+kMDY8KQrCVfmbKn4lz6lO7n+Cq8r7
wh4tKXjBOdRGNHFCFQpzF+A7HyMp9b2IuKSQsbgA9ghYd4HrXlVwl+4bcaW/d310gQSVw9EH0x7R
MKlHg3WLIvjRpag+Ff2GhlB0U08vEmE1eodprrvyQ68qpEpqxg1e6eJFWPHOUpjfgY1tdCsbYnJs
os1goBqYelXa3t//kQ/6Ac4AoWmGFNVNFOWuPNfTeMwvrinn1vPGtWdz3L1eDTI3KT86KXBk+FZo
hxa3w/bLQrBXt6iyWtcqZQtOOhLTBRdlsDHCpDCAFxrqt3I3oyrY/4H6Jgh9KSo4zxEj5Bwu5hYM
Oy1jw8MQ0gsI80DnW3x+lCWHae5ChQt8NcmbJzEiXse3VIt03rpKmuO2kpAiKjsV8VGyHouOxkVk
OLoNci5jgKm7zPnJVONa8AqUTG3CCxWK09WfJ0vKGK3oyHOm27FwI5kfnjWr+FhO1ETibYKOtGw3
JZc/4HsteZo+jI98Jr0FgaDEqs6v5uLr1Dx2ApeJXgL4/mIKI/sE/6vqjHEYq70iYMJQsxkg4kHT
xgGig73wt2sSxg+peCNCBPU25KvQmtOoN+eSkqQhsV4CbePPy0Cxlg9/ZLOiNWHaDi1Ts4Q/I7Zt
hXu/51TbMADrDRCyKXahBJcbYULrbU3oPenhP4B8bPPti5cvwufVI6SGHnIwZzmUncA0MHCzmoBv
f0mFBhGswhczeR7RVPVW/iVwjlc3FjNmIDu4jX205zPm/s+tnRxZjMtttg1UT1TqZdbE7Hx0ByM8
jTy5SKewJTVumcYtKiI+w0S4wtqskhjU5hpsmhUx9YWPFFEsodsM1uvinIlF+w+I8q9FIRni3BOC
pUVsixURwhlx2vWzeEkqYuAN1aLCqrtNXNCFRON6xC2p31VXFTqSzlJuD6mOsB4uddgohiyF1WAt
rQkTnNbErdahIfjsywA4SjIq4xm26NG8dWtwx0rK/QSSed7XdkI+1z7kHlGIwrXDC1E0KASQh7KM
AHAEhaO0NlCl1JnzaHgcPko/5SQv13yjQc8TupVif10137jUGaL7rDnv/Kn+P0jiDzjMIh2ZTWIk
dv120nPQnDycnI9GNPDdQ4Kx5zESGc/9vWMcn9DP+HOnT58c/XWK2w9FybZF3jQYJC7FGBt1LTS6
FuQHZPqxq4ewzLblzVNsfI5CUG/9/aNqvHndNtF23zIliUSR2EQRHZ7wVPxvcE7wmvXw5wXhhRcb
u0sDj4HA8x15FonrHhHscVmJFiBbbDc5r85hQuk2Wt/5dGxLNNToEe9jf9/84UlKy4X2R7O7JdfX
LxravwxoYAJNeVZYIPEY356TFxiGDGX6uUbGPhgawpSkDU9yxSUcVpv0GIm81MPAeN9ZJJUX1XgX
0VyZThpGLryAo2HWpegeCwSJU2FV2oVs8Y+3frHj3Tr+ZtLhz6B7pK+v8v70Pf0jA865Eem3YUF3
GYmBnjzXv5qh0kfR3q35WCVNRatQv6SZXb4hwNAGnXW37PAHiwVDiX0m2Yd+sWVnSofzX45xrfz5
atgLa0d5l19ry/J8pMBGAYDD0J6M4kvWmUWDJGNCATFpIDUgSXiTEXbV1cVJrNnL6oTEzAnqPuq4
B36t0E48VLz42OPO0wXyaXKVlxpH/+XCIO3jCHKN3TP/WZsvImXZbZ1qaon7B4fwNz87kqUl+Vuh
txZbhMQ/El/GcfcyjOurmyowhkESEU03EXjSXJgGCzif0sUj9QIZGON0Q4f9Q6PCE8meyFT3CWuK
lL0sq3UwadkQFue7TBbU7Fgw2pvrKW2kaeqn1vEUgmL3N7gdGgQKbT1Q9ynwvyCuQ+s/kJJQchMN
KwvFTpSt2jnkMZP7a+JxNDVgQrFFJpTMXsN3xwZIFjmNHT9w6QTfB0dVmHoxG38zVwn17GZypgyS
lmo7LW8Ifz7NccFcagPKF8z3RjJAZbVTj6P/v0xwhYa15nDAvLqLDRtQKPuOH+qskK795D4apGDS
hfjFyf8iyN+KaRCwzPYMSfl9OSkb0kaywZ8h7xplx1Zip7LmIRxoWlN8EFvakdbr13QZva6zEMdh
zzVuJQIS4ooUu9n6yqrFpSNR0Zr25Wf7yFnV3g0NCFz+hr0dOZWh+CwqR9mGMDY0KIC99XyZaAGN
jO2tthhaXf2UgHU+PVz070tkkDIqGknH++r1ex+WraPFb4oFQfJokQS2JgpoGpyCfnBdBfVBM1Yr
UOT4yXoVsedwcId/2GDRu9Np2aaVQdkuHVrXiqWlJVumzehUDzcerZtAA4MK/+8JdKfrROzOwyTT
eruw7+qOGUO9SAppbZRc4OpBDOe5F12y+d8y2NUuGbZ7fsspk5jnsO/XvfVcJK/y1ZWhAVrNfZwe
DA9kN3YgN0Aaatq3UA6dBrBqP/p0c8HYCY826ou/tmcqFpVEdRqU4tbrBTgzUpnZVvPiN6xJPqT9
4J01ZbpmkfLFZcBlCn26HtyQxC0v0eTrFeICnmSiJeQ81Ttzstz2wPOq2njbf/t63ttc1ieg735H
f8SK2T8FxuLRAlW5DaO+r+UAGkILrAHw3LSpff4h9lmDpZyGEpLMFXLQNLFM1QJbr/Bc0Tt8xYZO
vfFO3wQic9ld5yewys5AOgii9nLW1JY0sBV4PEa8VDuybvQrfKfiOK2cA1YxJdA4Q0YzOC68LXVV
3ACwQUF/aZhnNvypJICwotqC4hMljHod4YlONTF+iVk53V0ADGqFdvC94ZRFVAMBkuA53NXNrlyk
dfgCIzWgV/crlk2dM5s0MsM1s9GiZI1xWrrz76dBaWnhlFKs80T5BKGqMJMGHW4oRAcg57JHZOU7
uUFWdcJotXSSvAwonz+pmxcRL/J9yQ4A1mfAgUW64v+BkBNI8kZavN1x7t3qLCvZIaEG3bNgvcMV
sQBj5mTSlaEL3gNDxvanHx0RcNs08QZbFywyZyMCca5JbOf06LzFX77M2oSQp8nAbecwEovaq2hg
sgbkaWO35CvxhLGqySBNawFoam9T2dmOlQop2dn3uMQkwnPXQnb6dA9xGFYpBtBXPOTjksZ+mbIP
u+vBIrpQvhe//uTn6Wevam5OL1j5I057vNnmsSsaueXjsD966Rji2LleVxfDfYh8Ee9E1qWCZqkX
XgdpUhYyNQ8mGkqr2LU9++NADvWKOw/heq1S3C7qReNbxCHGJhdp3etzALjiB2V8do1hNGWeckA7
FdZsYaLBEZM4zejtt1fy6aJbblolqBCZ6MnlCdJ5ORjdklXW6FckwvaprI5nv6af3GD+aEUc1xyf
BEwyGdW2G1/4xq2rS5CW88CtDp1o2Gq8v4a7ifHp7azl5lAdKQGdgjCBu8R4A4RRVt4VsbxGxK/3
18REbKjwztxwNvJm9rktSMAwjiR0nm0vD5qmUpd+89BR992bEnD6A4ZAb74SJKiE2Alhl6SzgPBJ
uxneFJErTt8k4PgmCSSCgacfycelmoXIVj2qXcnMnnuM5vI2vmdCzFNwxyN0cBbnMQ3XnMtdI6J7
yQrIzxOVublNYO2fkZKFPu+Bw6WB2icHFZji2pqPj1SQ6dogXao94rYNvVHhHn3eSAWpDPMsEShG
AgGH4SLVJ1ElMrSPjy1KQkEKuR4of/TFJ2hEbKEReURDef00vBsGk6ptmNvBfN8EECzNW+bpvCqP
Nb7OUGdbyTjhpDTOM5IwzV1Yj4U6CbBugiUaadwg8z+lYvPDIt/Ef31hbnw9e4UDXG2dReWRLIJX
UK8zkim+2RcV1848Z1M1ywyAEICsMipwie4MLxz5U9VCE2C6OUHME1kmswGwJjeNs9PQn7Elot5K
D6al8/vNZA34Wst/TYl89CSf5JaMgLIdx8XLGk7RMGI1klLB2h2f13bTsWx1Hry06+cegKzk8Xei
JKl80g4eEeqBXhshjLD1/plUwTIAZLJGP+UTOAgRKk46jVMdaKnTk7CfPS2HC3CI4GrYP5vWNb1z
38ivnG7MY09afelnvn5qflSRPL571RpctlLhNbxKtGk/u/T9EqSa+s7anSQtyygy+a4oM8e40lfQ
NL6YGZhIVfyYrl6PzlPOeqyoEhe8UcGZ/EsJ2cytXDNtJ8HzsNAT/a2GbcZLME++kQblQXVmW32Z
5V2vPxuYObHUF2p/Z029UzeY8YrVxrw6MKbxIRPOpxbM4xIdlJm+ulsWX9uP6x6Gh3MYeyCyrzkp
bvFyeJXy+TaFb1jiR5YQvKPk9afQWXwERXJvhc+H2jMvX8PiwB5FGvG0wox3Vi0GbsWmxtLngOi3
4RHOsmjTo7VCJePLkzJmx7hLYDP5vDdhQLCCP461iKgxKdxdMhmPqxCX2kvvOLswtPx5w0XAWYVJ
KYLcKMCErLVQ/VByK5iTxzvpZx3SBh4DQd+4k91MK4SR9MV8llVPHk+1gIAvSu+NKqv5iWlotQnW
rErXOv1vvF2FTylHfo5QT6QRjenI1GZ2IJfAajbS4osuX8CPhaFMqm4AHkBiI8dqg04viEeg2zg7
0baaODFUimN4uqoSL8oUcRCr6jE9dzJ7s097jpTvnYTjRpcnXo75YAUI4P8lsdxeMF6SmM3fzA6e
Cymzvv0i8HJnsFZs3ivC6BAirNLu01huz+S3TkeW2k43HdNThyCZ8h5ZPjPwKbg003yEn3iWA3vz
e1obz8I0rNvnxPgIe7BIjKcDpAbp5rbQ9/BQud+yDdsMEpVC/k1FlXMm+BKYtB9T3ppZqeke3etY
VtDn9PRsdPuUhUy8q6mP4VVeuGbC4rWFfVE891+85w1OjOCtcHbjaIEe6PI2DYwPyvH29w7PvM1j
zyB6h9UHXJitGW4mtSnvQ+Thloxi//MVJ/q0AWawWzxgsVmdsFyefy2jKj18KEaS9nIppnbYFk2J
xYFYoVxx9Yt60pr/TFgrbrY6PB3bxElcbZ80vz73lgbbiZX8t/vAWrPdCohkJtDn261QqYA45B0S
6exAnx1n75lvl/YZJz0Bl3r9JPj4cjhfAqxJ9e4Z+/c/x2el15ZydoEYgKKfO4AJkhcxi/94cAdR
AnRYZdzPoh4eJhX84mNnAtu+QVwaFOj+Rp8MuKvNpTZjWqiutgQqQuKv7c9hY1PGahWbpyEJoUgC
bJxQX0IRxVB1tenjE65rq5T894j0z9e4bCx6n0mPuR1uLbbwvqgIeOT9/VZkWvJ0M2AEVmwc/KU0
jia3lGG4z60K8i9JJf7yciwke3uAQQV/aQBlfNSxvy2C+nTOnnCF0tQPi1uMhMtbid/CAS6WrRc0
nWZRXSEGiXJxOyaWyH1TlPCHt1zdgIxl3OidCJOZQFu+A205pWK2lTlR6snackYWljYltIZdqyIh
k2+b+fS5Fff3mrNWLkk3mg4QNYqtqXka9PqAOE74boYyaHNoM+WBluqnbTel99ujfaDm+h3zCSUp
KGOqVg/3bZKLq3RMVgEK1ICRAlnxPsnZ0IByUxXNj2hb3YczsIFW9WHkzXQWQVLv1UiQKEzp1xPf
N1xeSg3tbYXxMkLEsyysHdPm1dJckkZ8aRiRGM+pA46IZH9KNqdEmAFSFNYqrBFbS2Ixi+ChNCt8
YShCaKhQQFPz8CJUeT+1mQ4R8tuWBu4lD/scKtHKg7+VAgRaZx5fUky5IKsk1614qLZxfIxeqwgQ
7ALPkhUmJ1krsmQRumcmFjU4fuWYoNNYrMMPge0EBlUzQGC/ZV5F3ca1oiq8cgS0Wij0BpjflTcp
S2RSxPr/ZLKyx0xOwFIEo+wTD4pErZ1qmq4DVhM4UnNDR6ILJOUv/DfQwRwQyG70QbnCHMWycqLj
hDexZag9lV5b8eqZAObwXSdqD+ZDYiR3ai44qDpRZQfXs3aLtTqlZI282z1dNsU4b3Dshc3cDTuL
FSdYq9zVaK2mGHG62burzY7Gr40PulMMO81s1sSLdFU8pXhwQ66irt7COwnmct3KRqnEfiy1xqR5
VNKPrmsoURuXP9Uigx5n8UqgamnDtfg+u71UM+29fKmqTCGXMufHtXe/aF/3hvOQ24a3n0pSq9Ez
ZItI3YGXobLKpvhczzy/vqClXcBkTMMLtW09etVLWYAeX5gQkdV2W9A7ayFd/aHElia3AMAEreig
zyKsqHRWBqiOwkM2w45gV/Wo0hjJGsNiglt6KCJyuEMRFbMfqg2+XBrQcw+67Sek5rW0PuIC63R0
IvZ6mZ5pCtSoil4+7nUqaWT66LOHLK1b1tHTbLWBK7bvoI0WqIJWcri6wJZvyki7f41YD+t0fyCc
sdpTWYcEAo+W9WRgSVkutL/St2PKdQ/+fqHayGjyDSahkCqXmHAciTOTidhcbdcRchrBhzOR4kqN
yJYnm/QCFDEdnCgGUBk27snG4eG5rcWHaeKzT8IV1YMBf8wWhhIHZNqdT/OS3dwXJa+3IU0fI90o
/xcdJYL7BlwKCMOGJERoyRGqRZBM24ue9nPKcP9WVwOvQW6X0cXXqq0fiIfv0icKXxZF2KJvTkuY
V0KibKVOEqXKaueJ72yio80cAcUKboI8JO1cvWyPTwS+Smrcpv6bDE8QyROKR+1o9TxTJuosc8TT
O/ExPOmmvs9SobFW8jdens3BmGYmj2Df3N0TdLPegxWVS6Mdq0zixSV4SdE0fKwQO/Kg1PPHFZrS
gp477wD0ggiYciPWS1ErKakS+8LucPgPD8ES0r7Sr8wfUD9oOwGEejqWRcKHxq2GwH6ekqX+pHdy
kRmxbe95uD8WE0CQW2E65S3P++stWeqFTdh3nVaPT3eKOR0QaEICrjDbvud6V1BEXs9tLrIjyrF8
nM1BNh9K3G6HRWJ6msyroEnraBvoGGcicRE6USJHjXMvibPBx86WfkGA3KjK0Ecu58/Ct1+cIizA
5AjGJarDAYs4VZaK0/p2tlwxGhumW8V+T0mo9Ixkptbzr/x8oi5Baxb6zBPlYK8sSTnxvhpJY7vn
trn4G5tsbpdO6py7hZs4+uTh+dQrPTln72iaCxAr4anzcglROmFI97zHmCLyu9CD2Ne1PvzJzCTk
na0R0sbgwlFCNbUY2YAVOrLg7EpPGZy6P2RBzLz50RkfQiv/RMI2uKdcSX56pUQAI3y1Y483NiQy
zJsUEiUdLBS7NrWm6vIrDAHx/NQEnqnX2O3BiKHJl8IXaSIS67ljPL6H9AjL7lFe5wLAXhofQVF9
eSqlWT5UXzQMcXIwOTaRADmXoQ0CCG4oPwD7Y0yJgW5uX0a221Y1YtUE5bzczBzpT3aBM8yh/glH
l/HkS8yu0XjiS6KM/nVud4of9rbdc3ubDOgJZw1UhJQISvufDEKOdPtdhAb8sVUgrYdNFmZgWtxc
E3knfugPz6//qSKTGMC1p1NtJKBfonFlqV0hqNjO9n3Az9e0eZtSVMZEIJfFk9y2+rRLDyLI9/uV
pqUzvwRcvaJZiPmLXsF+7KzuyVWBE43cp7B+Q+28oqH45+sKFBrwFDrkwUuqGW/j4eH7oBb1CaTd
MxiGERVaRdLXyuGA2P5H/gKJiENEmJHsF/avguWEqQaOhvwaXAQUdjGfE+taji4jbqoepbozW22u
Nf79JjvGUw0dhZIFElw6CkNgwiDypZhePvKY+lvGmuYsVvHLD/Nrflx8aKVmSJ23znG/NQGrn5gK
oWeJSuFZeyHY98lL4V8bfyPDkwuq9F9gAf/weQ1HUxANZwXNuvWg+ZpLSzxdIMksrreNRBpph+wO
/Nf0Um3brJ3PljQ4dX+6cSVW44ya04GWfQC0zD5f1R5vN+Pe93ILtjTkfiG/p8y1QDjXmgDVm2AI
VsKZ1Mo6xi9zq949T9Pbn/3Zv60kMw0MY8nSK87wO0KdTLdYy5fNDGId3WVhQBWu48IoGYtujl28
u65jQRP58yeXeF9NGndL9PwYxYbArI8MUifnTLk+E5Jm++LF5xadPD+FvGCMSapmqI0x4+qatoGy
SkdtQIbFVF1qErxLnaGMWa7WxjPDILyFci6Cv87H7gZyrVMeo609FsJhHq2mPSHbkD7cRAj9X5M0
TguOYAaTfWvzepfrOWUW/xiVhA8/bBfSzkirl4cf2r/rmXOFJBcyI5KEIttccFqQZzPviM/IMdVs
5qaZu4rBJdkSne0alQ6gpyIAS8ZjjIXDs8CFF1Od7UFTsI7u6TdUajosFikZ2FA4v1f8LNfEZeON
ZfJziC8vtk9Lhnxv9gjVNxwtGJjBSyxodCWJLi4EPj4Zd9hZ7rzW6Hjcv6fglHcJ0hGEIDiFzR0Y
k69wqAGSDjX4hUHU1KYZmwnmXXFc/arV3cxxUx21ncPU/hLwSxJ+Bk+XZqkuNbOtzcF9jdSW5PKn
f6pUM2UFdTfCJfLcM4DU6uBv/1geBP6JJWLiQwtkVtupEzPfQ+2BzkRxDRiMhQc5ue0McNm0urjK
HEa+hBu6GXlyTJPJHFAcmrVSK/R6e7MtMH5Mq063BocjE3GayU1v1js3AUdWHH11zztophoB3eSy
BXg9SBQ8sToeOnmAoN2SI4L5Zf3K29b9BFegQclnWl5bO2rawHuDqN5dCRYdfXJHDQpLEAwyo7a7
/J/RDdJcf67jQbX0M4lD8JTY1ylqWBzj+K7ZGG5TDKNpNCXRjDIpgpeWOyT1jXRIF9Cm06e4tIjc
xg6/oB/BwKYn1QYDeE3OZUH52MpFKnvJkJIS2hkgC4Ygxl5o1uINVaJLccBOJFQeQyDzdJDCt4TT
CKCHik+aM1tKXMbCRa5JmIJjHl3/kOgr8kWhMNn4J2CBTcevywIH4AJ8wLTg8hoN1gmiz7rslStl
R5cDyTNQJPX3uBbId4xcUREmyT2K08r5ye2lghcUr3LC8OtFgdwNei0CbVxVJTPjkj2jovaIUWzS
/0KQRJMheiRcbaRWE9uXPvxbZodOwpjwBxOnsJ+dZZ+udE0PlXY8Y36TH2FSg1TVpUy+1XD7woRd
D9wQtOJlHxGzzMZ+7uvmXNBtstjDwtwD1UrYB9CSDEKx3pmOKC02esysq0Qr9bRwvAkpTBpn0BqM
LFHXPFhrgbgRwte3CrThx3wRVPwwpWdbVCnGsBNcft0A6INMMc260CzaIyw5S306SAtZNjXvTlzr
O2m5SJ3BoINEhYJmQc2IfS5rKkgQlH1YxID53DHQKL88fobphIvB1XvEAdIfy/4GvPdwLnOKsosV
81Ejs1/2S9dQAPBcBAlbKKCE7LlPu30f1fIH3qqIewuRVNKU+NWBKQSUYK9A1S22w2KTZR0CK3LK
OJsVJAMwGWIWcIWsp6Q5C+AYg8qWlUnNfz1R0bJOUAmBe+Nz1q7xSoJNwut93YGBJGLmGEyIHngR
fbSYYq/ahoW6573vkXy+nyhv+9eVmhkvPb1YBvAtbsbfFf1OuHkvzmArvS3NomrkxRt5dUmmGT7q
+5QX/G7/alx+dlc/SCHJLyhiAa57Sim62h7pwY1mgISkknCxCQMSlNDG6gKl+qItio/w1kUPFwru
x2WJERTY62JS/Two3Qn7Ez2C+B6e72ZaAXrRxumTGA332HappQY759yt2+yd9MzoBh5uOhTBDb04
hAZFGwk9k6eCzPIV24FpXneYfpi9agIKskYiCb6DJWq976OMOhILETXsGn7TBliQmiDNaGQGqkg7
9NN1elUA7LUE8jcfAz40VKWfe4Nv/NXcQ0SJQa3KbGwUI/sFwG4+mVjLYHwQlAxW7cFocRntOq7N
30TgAwNfne9amErwjq68CzQ1skh6+4HJBRmZvJDzPVHPGoA6MSLPPyeB/oQqz4djqHmIMOmEf+go
kylLv9j/I8NsWL89fzd5HqtVPQeEN/8oVThREDs9FchwH3CQP8BvJrIJMjWTXfM6rzNkCZto4eDc
TDA8wCBLvs52RRUhtCaPBxvsLCM3vMoI0oBr4wqJKmSEjsInmv+N4IaVKs9estsSArEs7OhyO7qb
ScJZHNoLGdgqouuzZ92vuDmG1IVU8Fs8leK1H5nSasjlZpVPl3ctjzLpqk4jvawbZj3Yezpr06yW
baFXjSHlK/7jMZwkYMvfymX/tY0sCZv3yGRDrGVaQXboJoRT88+wolhNIv7pn3mO3BJf2Ulxb7ld
wiuu4VexxXqqMUKaiZii7Z7Rhl9sGjyQV2JWkrfu6Kb5pui9sv/KsVcqTpzcJileYJwcV4bSD/b3
Wr2TxZBHkGbYPTi4RiQ1YpbzFeuO5YkOVOz538aYjn7M5kIFa8suNUPO5qsnjJzCQsRXxyLjEHzt
jCVVpZ9xP2FD/g5QEVy93WJRLxekH9IIIEiEzosIR1+r8zPwaCj72oOvskj8pDwzgLuB+VjZrOAq
X5uzkTRM/Rluz2UXUaFnpRf9NWaNCAWto1akiTDrK0eS4nB4mvgNdDtXfnqGb29IOszqoClbZtZs
f3zdn4st80d7ThvAE6Qpfet4Fs0Gf5Vyyemwxe9GX0P88jttM1FnXPjqYZjVf1jlW5jYp+sUVkM/
DwGHYHVHIjOZ58djGAlWzH4lNza+RlThuNXo1IpMK/tsyTphFOlLfSjDNP7bQSlogGGYuCoLFWB0
Z9wdd3LAdygyTF/4WihxvI3De00yV540DQgjFF6FvzWGQealTRPz+3nf2o31Ynq+F0NeUHZicMFo
jZErvMDC3Q0SvgFhIFo99ILj5bANJ9tFVfMcun7f/1N0p1m1EbgLhlbeJNlWWpDR/soawRd9Qbat
Xc380j8V9T4+U7C9EM9g4oH3SlQkoQ73EeS/M+bSlY9hx6OD002LhmZVy2oAAlB47Yy1ReiTHar/
WcZkQz7fUMNpmBByYVOTqMORkLY8555cXPGYbg5/rb4IN6i8Aw0ev9JttvgNIxPrAI/fO1z69y6D
1fId+TTxycxvREwzaUfNBob4usF6FzoHvoncv3kZ7DYplx/+TyI+dDgjS4k7QI/hXn19+xg+zJqe
3pof6Msr53lBl5G3OYwRhGO3b6Yu3sg9iei8m2QpPCKEsyx2XEoh9zHxrCJkxiv2TRbXQ4dIEmaC
UXoul9KQ9SNzCb/8swG0iHy6BCP7uKSVJRYe2g7uglRi2OSmSc6ZRqXtBfkCHy89bRkWK1c9lH82
UeIFGRfY72lrBvj0gE2unvqqUi5OFon2PLwWDXjXNqNR6Hy2mnj395WzuyhnyQD6yJ7601/rs0mv
T8IczjAgEySg4XTpqroza5TJF72/8AmKeJAmbPJSYTdQo/kM91K84ZqPk25l2isUnDv9WPjysFt2
6PddCMXQSNcgqKNcDBRDWekqOqD4Sc7cCjOKJSV2NehvolObYQ270o6UO0eO62DGM1hsgo0Ma+U2
q6sbqXT+xdhHupa1OKXq2Ad6i5r94sRyFLaOSZ8aerzV+Ez7urN42s7TjjZda09mlCxRD60qmvsB
w68EXxEu2Vqhaw732pzUraAt+rKbI4BXDOsKJBLeht15BtEmmE6S2vlL7ECRzPUD2ahn5FGyul1X
JGr7cmim654ulZB1QkkET0xQLrNg+2tS6ncQ/LcPjT4kOyZcVY4cH7eyIIOt3UiHC9oTZn5uTN2n
X9Am8Sz8QRdcws+T2SIM32Zhnv9kEU7Os7xvHNsNz9l5XbA9Xm03qrSU3lSLTYx6eB6z2/darm7o
beTrMeWKtCPv03BmOPtjZYpdAXM/jkn5OZW7iz/DL6EERCH9nkt4+DkQwRWUFAKwWs5zF6s7Z2fu
PFsUWXRtFkSFn0K0P+PH7NKhUzpU1Oj8+tgdteZYFxgGrMwlsMke/ECRkPkCF+0kEWH2DQ2Psih2
1egMCrfSMRAYLdCSruKGqb0LL+RDiMVcBGJtYWwKTn41rWja9vZ73w8tXXe7K+D7v/pEtgMfC5UC
uQqAd1OpvEZrSohUCviulzXmSfK19nUJEQikeuad+MXi+zTUcJ8nH6+ObtixdYrZn8oQqgXyM/9c
105hBeBakfkHoT/vEoFlVhN86ADik1dsFCVTf8H92SCzLkrDIjG1rAhFJBb72rutuffdaaEhJ+kl
hV6edNW/23f3DJ+SyzXgJVxI1BUXCvtRG3zT3xJK+tC/h5YHLwHaqwT99ol7YLlHbStYHlgxe+in
n0HjR4O29yUvH3eWEBtqGxHzW2GD5CxsnLEYUd5cbt5+ac6ZVWvboU/GuCzs1NfN7ewB7SNhJ4fl
V5Ty/MgPkNLG82SgdnApQmhzlhuKAmjkQfgnR+XN+yA3UPvjPhEWTShv2eaKV3qUSd4XwdL075zA
FYdiD/Io1R4SbB2evPv8tMwAgXH1SdxKMLxYJvUIQbIlZYwoVe8z2UWmgRLN9P6PynTJNHVzLe8T
HTvCwi3M5O6nLN0kGm+yi34E2VcVGaNQmm9HZITLrZnWix76aFko1qAWcHzCotAFhtTo6xzAjcOz
bHcpnrZAG7n8POOyPE8fr/gw7mL+Q20npWknyfh2axQUG4crutCSxtvuX7th8fFryDEXmtyxs8DP
vvWEE1/PhiCz6cEGD9VJzYLLgdAzCFfTVy4loHYt8vzoRDAuJ3AlJSPENUNznOU2haT1CcQA2iKF
zimf4IQXIxLq7VsNudW448Pn3/SQ9C3dkqp7Dtj5AIdbdtjrCGmyDuonKKjG6FzAauIKVMt0UZoB
iHRaE+h6JYtFdyOmdj0Zw5ecdpgKEu0u8LoaIvy3wOHX/ZKi87y5AnZEKrkQbHb2b+u96JAgyL7Q
EEY4VuIJGwqG5Qw1RpkVOr6767tGhMdDkisbzjsrZ3oRmGQ6i9lrkW7vnsbS4uOj82kLLWWtWXsj
sKqfn13qZjzCd9cfzwnZ3/fYoapUVISgdzoc4d/lYcxeoMVunzt8K1i1m5mjFZtte2jGSVg+Labm
YzvLKpPvrEfJ70o9IdkS6/PdyiO+Ay9Dr6CxmhBW2GCN9f6dCn6FtnxRpidVe5H1Uor9I4AHlObU
yhuT3KXzN+0elvWW5XzgUhYzIxjw6nXz+HZxJKr8+Zn1QO7/nwNPE+cTFJ6bVn469TnqYis+zcd1
CRi9rT2EFSiWoxFbGVR8GE+7BN+CWO8bUOOTCKoGwNPgdaUI4tSVn4V5siGUQbYt7jiszk0bGZRc
9wOLJwN9HhexEwSvzBHOXi4sQQ38t6MVlzbTSNGNmtuP5881OqIqY3Vqyv4aSLbil6s0tgqPfahf
3y6sh1yF+Y4jbkDmPZqkljUpznWhe9+Ru+dT0LH0eRBL3Sy1plr95dMzBaNvFcPlhIqOU7f20jNr
S12gstDJnzqsziveBv/XazwXRwp6m+LgybXyzpOTf6FPhofqQJHHAh27ZOSKkb9arT3TnMDEGRU7
TCgjK1DwXNb2K8ETyOH+9AagqMmouYlU7kw4UI6ZI+UCfeJrsxKk6oWZrPchevL3ixMhAIYaYFmo
WD0HppTvdAGJ+FgTOTIfkaBuKWhEoliK19mGDy8vzHUJlw37VJi4qDMrO9rLV9BCH8u460/oOaRv
YZERoH8SkjcsMoJdlIbXX2tHbqBVddruWecbIpwTar4py79k8HqFyB81PL1bI/dPzMLGX4NJRZcQ
7b+1hkJHKDMze+URRIYdJfYQZWE3o0fhhYGL7VBVCwQy+YRHt4RJxN1oUkC0Tn2TlR4hNdpKUTJX
HveEw5C2f0Ffvq15Gabwx7+vTPpxahYdT+9TAIsgg+60+Bupd4/wNCTMO+sAiSmOckbC8PriT9iZ
tJ9B0EG3ioF/0RMk5/OLMLOI8DMPzrNWp+aqTUn+v7v8JJdVOu/CpKMaDfoctZzJg4BTxhYY+2Ky
dzzz1y2qcGUHxDTCt7xVup0YHK9Q0RloiDLgG7n9XbXFJE/i5K9TMNqEBmeE8WsrK8daVHEVwmUE
ZH6kwRb+pJYoMkp/8V2lHGWcjI4SAAikJ2xp4rxLTPznwe4YX/PgH5V0p6fnYD0Sq6hIbdDrB7oI
pyD7N/BFSYt+cwjzJC3Z9c2x0ZIqaAEkux1FVUUmUtzYf1NVkwqJC5uXhUtUg9Wli/95lc0Afl/x
z0iBprjtZHK0yW02WTkIId22XpABBMaFdyOmSIzvLQODgDVzvBPlN9VE91QyflcUXjDMep/iY5cG
dXL5rK4b3phhDcpbc9noN6u4XpeBsP2Wuf9aO4g6h13q9koMCFldAMWtEyDKNx+qYPyIl7LNUgVB
MRn97WHD9fIgsJcUJvrfzGHOj4nWSIjB4wgkwZdIYxCZHYqFJMsbmr+UUafvUzGI0qo05W/ZeAPA
AEc0VkE1IAk5ubEXLQ7y6TGlbEXe2a9EolEf2Kyjo2C/wxTBeBLb8QxINavJWZbr66NRrjSbu24e
LUN1FM8eVbwpREeitnoLvEi6uUVX9Xsi3AYLWP8Cubc5J9/ecllZeme0M1+AfhXpbxqDKyVoJQBX
+UuaeU5m42AQs3gQPmkG6vPY4urOzI2nBoR1m6sCFil1BGxVCfnYoRJTibO+b/LAaeiFQHr24mFE
7VXxWZnHrvFHDuyIybmWSEzPcD7ZqnnO6VXRxWMowh1V+ePiwgixYcNjxNGdhxjSDiKc1LT7ikn6
qwD0WlJSBwkNg5+Kz3cG4GZWkmBuF/T2bDOwgyh1c4faIhvyY3Lgls2aT6kg84JEtIOt8Z20zF6A
hjJOJML66qAeeketwUiwK118LOExex2EdeSZbnKq13t1rDfciRNwywJXQu5VdmIgudzWfqKpE5wY
2SG0ReVD9HsHp5euLjANXvTAhsMFaGnELYtquhl9/nHkLJs1hdHwQLd93fYVftBPosgQb0CIE2pW
Li6WX3nrijgXIH/s1BGEWAP4XEBtbmTp46v27Eia+X/vD6PTPtbqDdjyg7NAbbGWGatnCJeDtQ0g
YSbhG9cVbQC+j8Rzh85KIH4gJ1Sbvyr859lsqj6nlvALlI1CAb11nfEujqDgwv/wnvK2kCmasCbA
0/ZcvudMu48rtXt7gHeA/WSyjGABl7Kt0mnGXI86fuym4P3+eaDTTqLl4G9I5Old3BDRKfUDcSFN
DMxIFwo2sAAsQAOIEucg3MQcRXTtFgvbAGVehoigno0LS9gVXP6LW8eYqjkcOn0q6J+IwDFSyG6+
qlEcJy6lvNQ8po7I1RkH0utZf2o/UFj13VY5Zz9SBepXOep8u50QiN56zPOScNZ3xeogWvVfWqmC
AaWBAeYU7I7xM6dAnqmzZK0njZpdOVEWrhqLfDxTrQoaHBSFiK/tFuDZ/LA4c4fQ4V/Q4XbhTKBX
OglTA6wcTYnGIaIjGtYHP4LFGnboA/Nuofr3YHvsAh0Ue6qqjQ+1sCzgWwrSIxnRctZAudOp3CJk
JzytOEY3zUuNZIEDYZ5ukMr4rko2Rx8YQd/hBqJOX7IcFj59CqUqA+0rt/MseR0TArX95qw28Vg/
M54RrDk7sRrR/7aDl6Mi+ahRM/OmSJSvtX5PZuDkhocYpiznCvOCOn8EXTZ+vKSyKz/QqV/b5j3M
YiGxeyQkSiWEcGmVUMwIz5+S5jsa6+3Br8MK+WrxEeKYbk6wvcl7yw2QDND2HUHe5KX4paWo4YOX
LoGiidpjNJDkdopDV1P5sWmMvbEP9RlZru3+S0Td2+p2ma36RblQjmSL+fVaUXGfh8WxRqp8GyFG
+8hzocuJxMZEm4K+dkHHYoaHhp1VSSCq632TvXyX1b11gTme/CzPUl1mD1Z389A/QEGptqTDPUOZ
4mAJIA5P0SkfiQYH7rf2l0dkenRwNf1ggLYK9ftDqGZREbRZSiAHsrNiST6r+AsiaE8uVB+pepFM
i1JIdVGG60vsrVVdJZf6Evffc8NwvBU9NrvHetzpAh4+YSCr243n5NOGo/xczvXPzEG8EV8FSY5X
sSNKu9bJ1PaaOf5+QC3MqQ3TB1JupWS1CZyhDzQkk4X0GsBREDAukFJ3kVKVlsFwkZk2e19k7sAw
BSw8Kg41FjpAz8ZigGFvP0Ktec8dZTdnEwvrOGQ9bMOpmXcAeDSpnjxTAtUhAw5EQ8g60qEFZvvy
36sxT7VWzOee/skIAKomE8lOd67m1WmKPNUQa0/6ytgbQ2hHROPz1zr9c6m1ns8/Y3PC1Vzta3gu
hSroXDUgUi+SVTvy/uaThKw4pmz+2vxrFoAEY/Ol4NRct0bLOdawq7iRnGytdfQHVe4NDpecwHg6
gd6UeKZHgxHayj54JBScUgk2uZEE3Cys2ZWDYohIkVIshWo9O8oD9uv+rF0+dLJTtwCF5JlvQhf2
reorWGsMOyC00CK8IDtof0x4vgm5tSHQQNeqm5pCAHhqcnXFy2qpyThJBRsF7dAMNbTJs5jn+h/g
SxoNRnVvOCHkWegm1uCQpVjx1dEkOReSqdxUDo6uRdMhZpDqo7fVVeETeMcuQzHubQ8HehqwJqUz
kq1axGKn1vAqCyFC7Ps27uL2zKwuawVu3MkxSUdUe5OWspVwdn3XJD5t5aIzBkORpQ3mjCUl0L9f
vNEmpZjF6tnfKMZmDOQ6cvOU5br97WAX6BqwEfGxt97ysuIcrPv/IKbp6NMhMCY2hkMAv4KJLbX4
6HNdKZqZHuu7h8651M50LTottqNhMLt/PWuSvvSUcuucmIFD7+wLgLFMm2hI3EZrm2/oylyCSvCP
hnpzxaddjHc0SvmeYGVAOtQOLSFt9RpoCzGINUJTBVhTLE8+YwxT8seLxJfPFxoeq19teD1xSoFx
x3uDePTTlxGrNqJkHymC0NM5jiN2EuhNIQYkvCqiuuMxmasjvGeKvaiQJHX96r1VQsG/6h6bgtH6
tp8D+Nh6WiHVYa19RbNcl+D3Cmb2bkH9ygKjRIUccVjtFNm53aetgkcdgUWJlz72E4IT5DpH4oXZ
yd2ymIoIRP9XodX9vOy6F/2k8JpG51YZyAxklqK5H/xfvnKwvmSf26CF6o1OKgEF41MmuNiPmbma
YircmRmFKi13czC0jQCvBGcsxYJ2aNId4509tTwnxsMzEom02ukCPluyZNRqCt6ikiQ2ToEqXy7g
yK8aGmLeel6JRLP7ZzfUxhQo8sUIJ4nwG/MPUpK55BWPUtTY53E3cXw+RtbUgqLgmIbqIgaOJLH0
IYg/vksEJIEG2ZAhLj9/Y3DSQIKLRagv3xb+smigVDIXKMm9/5eZmVF/Mj8BG7s5WQ+P7KO77XZz
59jm2zjfE5sWmd7lbP1DjwiRTsbPh5hBUIYxfxLQNTo7JhMUBga6KKWwc1H3JHw+DWB0LtKFSq/Z
BuXjYOFnwSGnDG/4NmolI/1longLg3NtFgogZgGGtG3Oipz4VR3iKnMo2/PbHX5C67oWATTsZEkn
Y338MW/hk4OcYsxdwCIAuKC1z1zby/tN13URfDqRJ6uLVtl1GX/cIin+N3Xu+2+w30Xx1B+5HMt7
Cq6U8EQzYBWGFEH6uJXGARXFhDZT6DK1090ZtIy1klRVwtFcu5NbmWV5knZioozmQmTw+6vw8mEo
kxI06JW5BDiHWirlYdBL01WfBnbCLeOdkcfbl9FXbTy4vIOpGRH/Q+P8xD7PGSqL81dy1LNdO76p
S8zpcPzcSQ0wUAq/yRcT05vObHb6yoor8LgTXzFB9jFvYNzMucfpNAl8iZMQWWxRkPoDMzEEb/DE
PqVO5MNeg82CLsTbEB9RJsVtxjhzQd0A30GE8JqQ/dyiRu6I4JdQlnTCyV4IHJx51vSZKH11Un7p
pxNGExfORDlgGcySYlecogTwzB6NNtqpMUQwfDfI/w1c3zeT0EmMH/VET3MhDXRyPBgO0stV36bs
lFLhxC33TuYJ5nrIGtK7QrCf4z6f/1wJQZnCO8YH6ps2a5APhzOXWnj/XseJdqAZTwYEwRwrg6f2
ycxamgryxLcUqp4q5tOedDZhHGWRfKMppPacXU83e5zqlKlXROySRPvGAbAwYljjyz2GynHYvdlm
s8zVbQpdIpsMWUJW+jnbQy50Yq9qKORsW8BJ8C2Vy7vZfPWrH6Z+kJAzG4W9VWc7grhlCIuLVfOB
lpj8Xq5vCVZ3bvgwjfJPjXAW6GROO3lR7kvWsB2M6Tql5+jeodp1E/l+vGcDCJKvhim1kjvJyUqU
/lkv/dSbLl0KVzeLjVgff7EU5Ssof9Onn+U29BIJvE50oHUBT0i/pTCz5b0YLm6GqCpPyPbUwEbv
KD+ZHdYE4mhKYDszRK/7WJIwHJqmqFxFm3ERu49r8zRv0cYRoRt9OvL1xvRZfUESv5g5dMfGP3KI
iWSbR8j14UndwdKc+bCIpepBq3IgwufotB1DpvS0sifHQuVrXV4TKUXFQXUUb7CewaNZ4kIyZ8bt
vDKAgyJZ50r2J9tp3J8xOJgIH3qd2t9JD2/bml/WSDjkZvJnZP6tp/ag6ljMGTZ0/5amgR7vzmbK
Dcz2lkFfzy0Ht7o92L4/qCqT2gqLaQJ72Wlv0AItZa8j4GNg0ec+CrCV2iiML8Lyyu5GoCDcc6+U
M9GeCbNEHA15qaqNk+1qV/cA0zgM0czdMZUjae5x4f9mhb11mAx0hZOoH81GugavH1Zcb7toleAy
BzFU035LCpDoPbNAwGcIBx5INJyELd5IXRT5baN3SkWC0QnAESOa3vffy1mKoZ+9ilggezyZs1tK
h230lqmQRsNf+CuAMOfr4YUhFfvX9LVG5gH8XlNENXH6BDUo9F96IhS6B7O7FZR57Y49rf5rbtwn
yJuyJwBv4Jh1CTXIiwgZui+NLj0R3mt93nP9/GBOkjZLORp1u8i+AU7IdjwjcfQItK+gmbA/qYNA
QkzQl65We24N3TCFE9N0yqx8a8E9cNDbzJLUEtqgtz49Qxx6OZyQqDOhkULVwr6iG8MXfUhLc/2F
dJrAgKm+iy+kiGnUNpFKCWU1hkGHBY3NppHqEYsr6t14vmIRJHA+4QIX2NRU1qMUJSSvJ6Khybdh
dKeeSxNuL06jL3K/gFJBQoH/TfqGzF/aQTpLZ/NUqh85tt2HavBWCikeh2ZonzM2c+HQwBQqgD1o
ZHQdRZmYUjVwqypS3M5nsRZk948/HwyJi5iYMGLmK/Q1vet3k5ClFRUlAdZ8LVL7FgDoCV6dYSqt
7ldEWxKjnIEfEPtM1sFDkamkJEEoNOV7NbyK5ozNqAW3/4VDMQJ8PFj+9An4GLIkoL8CXbtFHUuv
sQY42DxamiBSX5rrbwiXqdyCu1CDtMOOKRwCT+Mu2KBaaqQhbqa147X/Xk7FihmKkIjYEPEJ40u4
MzAGRp+YRzH2fYKcPiJYEUW3KDdQFvynNpuRcfYnzOMHHtmv+Jsyab/CcaS+mq+1KcjL35GdXH7g
tzl0l6iWaD7HHtpUDPOjS8TV/HNNNoNupYMBJqfXStQXYANZPsYj21KVoy1CTS9TGCsFs0UAZFZb
fDgyogtwzybcOilhfC+0reYhmmUaiO5CkPcymOJuCfXpUMUtdP2CmK1lz0XhGkL3w+ur4IMfD53w
SAKim9/Dn/4WB18sZt3WqR+/fg/sHoPScLczAW+p6Fb2IiK3dAPHKHdh57V1bOtbZ7U79gpK0GLt
ggi0Ko75hrH0bl6ls7CW/R+mLyE4akmIogNLBTJ0kWNdR680YDl/zcpx55M6G8BOfTKdoMKEPAAh
4JZfUGrjFmSW7iADiGSB27CmDZ9SlyeS8bAbJ7M7ua7d4nyMAZawh72RNuDXsEefloJU/5KvNU6f
e0ho7koiJugPw44ppuA7BAM9Y1UeSdiTcu8xMPw6hJadyX7ubKg3miLteE/J1sKml7nKnNqah8lP
jAHXQoTtMeml+4rbEXLoFflaYIjlbWT0490HhJM3ZLBGfgz/6mTDiHxZrqQqX9ALwSqY+Fgv5mLc
HVnH4FRONZUF9XHO7KQ/GF1H9znpz00CxRLnUJiQDy1/58ZtYx/ghAUmxJ9mVrxwV7Ia4QPxFUlV
TG9RhnoRuo8BrzOagC3a8bqc3qfR4Gm007Rmn58luKzOfC3+urd/oPeKDkZEAyxIH1cIzQpaVWSC
rsAdCdxEolKMwfk9NIJRMvONvXdL83l5iQZdOuyLId4RRjrrjdPv/Dn+QLDwTIoG+Aa0NGcCzkcL
10taY/sH+n/6IR59FpRx/VnU8wwTEaQiREvK1Iu8ZmneIiE0M3Rz9RwT8DajwtRbXe9NiTol7Td+
2FFGlAu0CKUGiQNG6YBr0y4YW9gIitbw/E3qTpaZy1gzBnzE9872eFqL+eVhii4d3d/kQ5u9Panq
R2Hzb5KvwYZI0F/R1Yn2TIDGHhQJf3W9pu3lukw6JuYyo9Qbs+sG61oHVFV48KuUkymV3iN1j81Y
WZ/tPyo3JuBt+lo3LFwYQhCrI3WTxUz07JQusbsKgjD1Lsg3vFQosolwXNHLKhAAfS9jeWgPMIZl
WyvHiZSJtbY1dEybaFegihnS7hvjjueZUluFwGUcnLIXhZeBVEmEYgp8PpJkjTq00sZKiREuyVCH
BLVukuYNwWTxh8Go4K8uTJeXMpCAIYjCwaN2jEZaHOXFPi6AY+uEeMU+P3Q6hucq4GLwWo9c/A14
xyzdSHz8LWdfb4dC6+IoSN9osoF+vGYdDvvRohODCtg+Wz4urzhb5Ex2VifYudgtaW7aouPoECtX
B/FiV36/2Ums25szoPLgLEdfIkukNUDyy8jFX1S/gKS8BCK99FAA18npcBwR9BNBcMmjXcumIgPi
RRtEvQa+nlu1t1QZcaOJQi4Szkc8PDfAQ4zeuLAAfRE2vc60yga0OhnD22TRTG4BwjfJjJmDiHTx
LYNgkdZdnBLnCJ27xtm8tew9DmnZIaeK8OuWOMLzC3tmbamWyVRSk3nyCKst+RadZmAxQ3+fP/1B
bIz9m/JWpWEm430jHx5s0OpfOK0ICGrRQhfCALc6uPhu7BcahiDT2d4a7eC9kFoRgthS9YSu2mb+
7IWo+QSj6FQNnfj/CYigyTl0mki1kaShQjok5J+3M264XDgMiCTOfw4Fb758pPIWgiNMWo2gbHec
gw45SajAOLdNIE4GqxFBRr7eo6ZgMbVByK1XsXjKGHJr0GccCaDs6ATTVMi/LwqUJDz0FB13Zgkt
XSMhWpwh+QuuSmkKOFJAZbCjks1VJl1utllFwo5Ifj0n/xmzVc3Rx2S02pzKXrfFYplmr6l0w588
uv4nSkUxR3GPJw0HZL+mJ6xGiR2F6ygS2ifoayIklY0VquoQ3qtI2DzJC1cKNgws2EY10Hr8Pp4c
68iKZNDXkwWN/8ldwTJjr1y5lpUx1V/wr+DJ5f3xHXVNir3ukegrgXVwkYThX36HVGys0ba86v2G
qGUdqkvLHwTF4LDNCVXPl2AJpVj1e6F+4xmNRlktoRH/RlbHvSP1FjcITaWZfWA9kNXlwkPcNcJ0
d1QG7x75+u/FX4Geir07KC+48RcNJrsTc/bWQ7WX5G8yb1YS1YUmRJ7F/nXavhoy1n+QBgCeeog+
mvuoZ3bkX5fBC4Li74YIKhh6wtscYYJwevGAREvvaqcFu6Qq8ZvKeyhl2kqeMuhi8Yjz2KJajNqq
oqCt6oPIuVblkUJrgW0WT3/WoKQgaxl5Mgv6uvleGuXytARI7fo1jdmAaH5UIu9Vet9qNeAkth6s
Dkl6UjtU9SUZ9PGRZvZNgegaumiLBPNKRsKUUP5Z59FPI777IfoCZ7XqKS7CRk3S/F2U8nrsj6pk
aV1p9/57kzNjHQBpl1dZku8YpC9EL4MwMO6O7L9jI7MyskFu5je9y/qYq6EADD3jgjwIVbMaUrSH
aPvMFlFJnynru20vieMdk+MuNy9Lc3RSnJshx9xDARqQrnlyt6iwJz/OafaMWq3f8hev+ULs+6IG
rGypO21/uLrDO5vylB1qrqt54EK/3eKre1acAlmZJSIYFbRSmti51We9mk8JL5jJcb3+Eqm/UL4v
Sfk5x1+O6zciGLWgQbDZK9chiZFF+UHaCm772f1pFqdETNarfn5PedIx62OA4j/8Q+zGdvpWVJFE
zX+PnEdODGM/lgMLBtyZEW02RlhPyOKnR/MKn0y74JGDJFccAIrHm9xcIBafz0tCWMEc9nNXucEG
Zc0/sBnWIILs+3i6YCkhgxA9p/PNrpvh5s2D2iQa9zvPTATRWSk/ijm+/kNq9oIqKue9yHX/kk4z
Aphb/okfNtOgvYHW1yMhQhliHYYfXiMz/DlL2Ll9wM4wzawYe8SLzFlV/avY16YCD1wF1qEyvoMu
Q7JcTteeRRv/bQkgjYch4dPEpQn4BDLRlkwf+ow0FkRMN7Jlsp0Uy+hLmEQM/396t1cCfnmG93tD
dqslE1pOiVcHV2PtUa2aFdqqhyuk85yOwK32XwvVOyExGKQGqSEmgl3TeGeLk1kpAsVpuQqxBZ41
H/ZAXVoKLCxvkbWTeNFCeWJzH/CDZL0rsWwW4ha6Ew77Ds7s7U8WAXZj9vcAW6a4cvqJnbxf4Kh7
aIPRbyu/F9IbbZCGGRDuYMxW0gk7ZoaWYqBilPx4OmflcjpvLXOknek4/KDFLfJAXUTsPkut4VxA
Sd/FfYbu2m99WP4u4r6L9cETKCjS1RKWWse1VO2lqomsYIm6tK36HQY85qTSzf1ibuoOAYjZ3L30
d7L3jKFOUL5Y4XpznSAgEt/9PKpbz55pn9JqQHJkPxVUry/oGpjsI7BXkXxaaKhlLkPWlFcpqYl4
zlzmBr1HNNmVsmdOsQTFz37Q/xgLaXBmFf4EJ7Y2q+5TUB09/r8ON0b8Te65JTfRfboKMICC7oCl
ULUqh8cuFPlwPi3kpEzHXbEgBaImt9D4E8lmtSqR9qfBPdUjDuf51frIIKft6TLcvSmOhint5fZO
tkZ4IAYvliL42428ohk7eD8VVPI25DBzhd190utbyvsDVlmTTM0iV+B2t0P261jZvBk0xugplc7i
GW/KZ+31uW9BQ6tGwE+CPTfc4FSpeXHUTzZ7N8/IZmAKzag9qVtFj/x8FftCpjRI8Azygoe8cYfV
pBeGeJN8CiOnUkWLrRQdy50zg5DCkcY5pYJ/khUw4deH5FVlEzEXQ394gCssU9w8OZXeOroXQsJc
QCgJu+HNlDY5qb21jaCOyJ+Q662qVu2jZt3d+df7lW9C665MIJXKvga9Hep1NLxR4o/IJadRk1V7
oYQo08L3r6DXPOg1LbeI9eDWjfzu+GUzEByFUIev6lZvkbdB7/Z4648y8q3/cFS6TaxqV3v7GK7Z
U/MNL5jEnvb8FE8yc2bSxRgzvfZqrA6bkcnZBcLRYfqAcjD63vsqMoOxRkByQC4vsDNwnxoIpTBZ
5nq4TrdTh4I/S6SEHjo6rjE8rly0PjOYId0Lab/oSkfZrQfl/9tnO+ULoslzMscRQocTd3Oc6VEw
e4YjtHQyNsJ5DUObVTvKGWZ++595flCCwBZfXhtnLV6YBNj3OtQwf7ex9hu64iz0BnoamNWrjhta
PjATGFUAcW/Lc9i0zbOGWJc/n5SHOJo7HJJMxz07LhGTWUX0vbOLbndX3kAkvkLV3Iubk0VW9GM0
RrGjvjE2R5djymC9QQR+6dnMlQ5+aqSRuLQCMnLQSRKbxY4b8kSVidR4GB18kFjqoWuCNAupvy1j
2GdUeI9HZoFF05ZyHC2qbI5K0VOkuZKd+dfZBBNv/iMX0SsRBRD0Dt3OqViKJZbi+SXZDK91iUKd
y1Hdh2iXqeCJWSKJJp9Qvfaqt/PUlYLGtnFSV9xJzOuO2oB8ZvhDgmWzoIVCgwCGxOum5+fowJHv
ZVUa/caBNCQCVtWIAvw3xLiVIpMtxzGa8rD6SpWO9OSHGOLsIJcbcKweCZ6fGNjWXlClRgILCf1w
S7Riy0qZElzls23t88By4LFLRVCJa4EY9n/VMKDBKrgU+JtzK4R3ZG1YQCQRIjD8ZU8LIy+HmiLg
JSZXCLqYvZz/EoGy4SQ0SSOarq3B2xVEraS9rbTGtizUhUF4wxfQmp1XW+G1eJDmXe7Jj7pqzzrH
16ZHf7lhjRSsxkQLVMC79k1H7dQ3Jy7GO5b3BhyDouSaoNbSB+HFLrSpV7TuRqEXloSqBcMc/MaC
CrZCxZj/SndT78geJVgfo/S4sac+YUB42fjf7pz9iR+x6duOurF1a4lNV9THsWzHWoanMTgQ/z1r
zq2yDqG+Ink/9i6UTg4RvUZh4d4JdAk5s5uxXHEIRFHk+/U6i0AZkEMBjuFzkqbWOqbuOf1UOvJH
Ws2pXP2MsKOhEUGzUrau/MMGu4s1pkXnzTwmk0R9mnLJpIxBkql1eTtnVLL2aip0eUFRHX8PnoXQ
PeJP67bklZg76efJQK18xpDP1OFOfgWG3IWOQI4Mw/K6e6J2kT2Lb49FrBxypZRHkevmnXgb+zcS
YPWcZPryfAp8891B1pfqL6rd0EADfN3eDwrqgLxFcNqVikjsTZfJURsL1rbUpj2SQt11aPKpy8oX
xwpCDeLHxnDhUZC7D66I9vZegWJsNbiu6hCqWALG894psEodeeZuLr9v89ECbE7kFp3EiRPafrYu
NX6Ncq42RQQlnBfwFDiBMDPIFiRl07SXoPdq+/ZQkUj3m01Dcumt3itQpwp2+IbstL6930cmdOGw
8b68P2mr3FxgIUI+QMi5+bz2zYfRC85luC9QOO6CpfYE/Cl6gZQP0yHfxWxpBG7/KtY5SqGMoFrf
ANUdfTsBEbLVQgS0y97FxeQ0/tSD6eYAU2B2t5dQCwGlxyrrzgNCln5DQ5lVwcoFumN2+W5bXOtO
c2aG4b4ssA/N6Wv/s+80UG9hMrnnhv7+pJLAafIRxrRTFTkE85Dxecc51BW5zbKUXg6P9y6f5Pk0
7aFDPWc2YjyF26QKjMEBGBNEQVZXfy8++GWvszFi7wRvEC1/a2r/fdcurcwcOF7WXJVTx3rD6ITj
IGv/pT/i8WFPjm5cw5Hmxtbp/f0L0VteCJIz+lnyWEwM5QMdBsez1AGsIOGVJ1wGD0oDjdk+67bp
/Y0nhMA+QCFROuzGHVfVnFruzDilBEv46WklLc7m+P/TcAuSfm9zsC5YKVmFhaQuprBqTkxLFeHA
g+jjjv/a5mwGjihN4tSZSDRg6/+4g2UYeh+khkiOrUcX0PMxx6usUZxUdh8XuurdbgXQL/TWAM8R
9ONtUTB2BjaGUSQ8Uz0qZskb+rTcQcfseUds5mEECLIWuejl4WFWyZbtjpNC4ujE9TZEDUYrFT/X
dC2PsgUKhGxu+ii+GLTG0MU0dIk3mFKKXl4YURYwpQMab25MsulqhegPTNZtOonrH9D6T8+RXXpa
C37/20oTsapwZOHq6l60lava6Ni6ACCu09IyHLLrqaFGQV9+AvEUKqOBUuzoKuaaNalek6CTpuec
aSjKRMPNhyOIsqOYErNaOLGCnwTVKoI8pZCQm1Ux1fLEElKRSL1hWL6OfbeWLbcaxoeCuh10g9u0
CfWkosD56XE1cRa7DOGLkHj7dr2kpanlD6fG3L0Ei+BJ9PvkbK8RZJerlgvGwwH3MOQM743gA1ab
ecDkdWOLyqWJ+gkDYBEq27olTp1BZF783BIL0GkmYk/YbcksPLanu22M2By3ihnJjMhRdaxfEWNu
N+bMPw6sG0HHT+uxxok/irdFNugwVHEVjsgqZ+i/6YkIH0ZJa1teTMNLtEh5sswIWRml9abDDF4l
Yll52jNdM++EU6a4sFpVAM7VFkAX9hHR7vlKe3vy4DxZ6ZbhDWHmMOzNOLl0KlfDsZLpQmMFH4CA
6aKZhMjax7bpuvWR3PrXe4vP3/mdnLO8IEpb4BE/rOoAFIIHMur/g+hH4JmIKl1ltPgtRUwjXYug
XKA5A+/w13C9I3WMjGp6XSeL773dw2GHhvT/NsjCemNOYwi8VoH9IRt6pUst6EdxU1bNDQjual3g
YeR1/9dwuxFygThwBcny3Rz+gn8cMXq8Xsj9dH6Nv4kMw92TayyXsAc45qBii2Tie3W24GQTHG0h
L3fWrwJChpRc/IjLuXXxxqSlX+hmNxP3nOhmMXy9QyibzC4PriYprzKezNhMz6RrSyQboA3u6fA/
XlnG8kYf9ZsRUuZymyeNL7ENotNmNej9eq/6TXh0gFtOEuj85ii1fSMmObtHzUVSZiUJWpafcZ7b
y5v74jnnByILDap4gy+FfxgVhPPxd5+X53iR5BbG4JWQTBo654bcYioRTzkNiFr7mnl0BA42fs2U
fw5OwJtGZ8n4b3zZAx8PbDIAO9q6NT2jZDr55AzppUgI8wbhDLujKkS4LRFJ9IRileOGkifMQ8fm
si+JF1btye9/Lzbej3nnNRvyNRfU7DKnjbtEXhvr2qfLc5r0hEJoPoHXN0T+jZvI4JA79SsYFDMJ
+hbvNgi8Ds335sCYNtU6z4aRcafH6QZyT93MWGk0+8JNBx4WxTNUSi8S0jQnqt5s9x9yX2bluR0w
aCh5fIUBWme+GZuepI3Q/18GItcz4ufsK7JADZ4Np7JKoTl7PLPqn5gAl32zr4vCC6q3AnDK8mob
vSsU40QbKPKBoLrHqVfmFwcYqrl8n8IH8lWfHOoFgjEN/IQp2IncC6ofeuZsywk94RQsqXU7uk4T
Kdhksi04km27TSecKRTbULjG62Q6ggqyg3gMxGZ2oWDbs/q70DC943OpQ4HyH8v5RO09XmRJ2T5y
eXBUUERd5VxtppXNWQ4T3WjjTh7FMkzNQDLRgKMQqJEPopcCBR9L5HKSx4rGJVCUGzI+pF7DMItF
XaKrSGDMWTBdCrRcHIEsYr+dsfrWgagNJlQcu/J2s+yD6DYgSts1ZeaUOn46prOrntbejQAHx1xv
Qr5Sp3MgZnlSSWI468mEORv8QGwCm/JXA13bUC4ea4UfmW9tEzmWKzKQ9za5AihW+AMkfwGAW7yR
+N2wxGHv9Gtbc+kJ87tmLffIUorHq5KVVgGcnjw15GT6Vz6fagyXHkhTzdjUPv94D2dNmgv0NQWU
PxaxwWMR+FMcInWu4e8RZTgCzFZBTCL4L8UeDBRVo+ChvOfy6Hp522a7RY+rHrX1eKDlSSMr86wk
fbnmT2e4hhmCzmksjF60u0aRNZlPSAbia6k5R1BtV7lUmzrWqF8lRxLFZrj5kDkt7cxcwkmS2/nB
x4BYtOzIgRb3bvDYY4PObSE64OryDSDtBxrGeMDVEcZ/8QNPtKRV6Ttk1EKa4KKQvmVtBSZZ37gP
DC7+3bW1qCVxGyX8MUQ3kg59sqQNKCvP28rQvWDwLsKoUIEKNFizzKJR6G8ZLJrBP2eiqHbqdC9M
Zk5nhRT60RE+0INhcg7YwJYL14lR//WpWnu3qD55MY0ZIt5yYiYfjV+/YOD0JrP1zhVTZZVfQ/1y
p0AgTRxi7A22azwYadL8al3squBHrSddZFYFGH0jCpjwmEuiQH7zv8o5bawm/PSZKtZRJq8wMywC
N8VrKNuSIM/9kKTRy9otg3s79jQqE1lyr//RF/Ggkb1rFNSaDWhyucNSx2WsLtycigSt7Ovo83jC
hG4Tv/pbYylYb7iPEJ61tKBV0ifnTgsqyKbg7e9zBOEKFjPUZkSAYQ1JOUaYU9AUcM+jvDn+fRWl
YGdmjt12pSSeqPBGClmAXeC+KBLfbqS94JWWQCq3Mh8erIcCeYk5t51MGccL5+wcdjtC8JG+wy3z
Q8PEqoWesdQlw2aPtiXVxspHh3gHfOBatJtSGADwA4bZEt326D8uAkjRKNiX+idPULQGgDrRMIyv
8MbRbwB5uQZBbBRBWiBZSsARWaMj6kqio9urZStASyYElv+GEv3T5lh7F1IMc2FGO2s7uw2IS1rJ
iDMh2tgAWIYkTIqsKmzUhLNCS97ZnP0nyyNBMEdCTW8d6FHssZaQo9P5/pgNoprItI2Nd28u3bws
FTz2dnnSxWAsouAD8hoE9XOeCxuSjZFbBjeMjgEaAELn5Ba/YEvMkMrkzY4ozEVEQ9ei61c9ubiX
Dq+nVteIPX9aSOSUwbqejfOyh5bwLsKFJRWoP/ejdOFGaJyMlXU1rSsd8HBTjTeyOUC9Al02odln
ZNJx2PF1hFtptYYC6Hg0Ay/qVRwgcjKp+UZbEe8lnr0MyauHD1gM+SJ9zIF9EpC4sPoIRsPQ/Ih7
+W7cthogiidNuCDG/DL8jOYVgKSjWfdxC1hsLiXWBOUqA9Dyi24+TLSRYW1YADTsopz2rwYDro51
4A0cWXGF1F8Tp5LPYMZGTB1JPfeYz7BY8yRuvShkUd1mJ6opA0RJy3f9YO2mti8eWdbnZi8sGphf
ULC4+kSEet0/w91RknY4Os029R+p/nJ9dXP2zf3Caldm04evEefs9AOJv4U21vJX70kiGykSn6bS
JXwYFzwcZ9viNzucGYwGYUON4bYpVtqqfYA8ZxhXcuOklbiE6GXQFKSb3PmxjKFNB1j0xnj5PUoK
wDCQImW5rq0TBOO71xRtDwQrnw1j9C6tUGT7yIX8pzwaLb+JiqSYKCFPUkTdCiZgTHbWm3SJORtd
e5fDhEvQPwdmtk4lIX7jp1IsmPFYcZM4l/xtS/zhe4hbYvxC9oz2sMORjczUNGPBU4D1jWYEkOCc
yjA+6wLdC4+PdPy8bjdDbTaV/arDC7NTgSIJOTTLOumqRl/cKgrkwEAGkue77YHXONi0CyybPo9g
15/q5SD7AHyYcyjQmrNaB3RJCnFWK4fcRM/AD/IBtkSer3DqBlNldnl62JEVWKiuS6JI/osJb+8q
cFVh0CUzNQRieHUk4YM2vpDWp+2r5E242CxXT0WNmC4Dk2kWjyluBmCF4Q0ittdFqiAivYkMskDe
5vSbTcns2RYJjY7LmNlN4VZXrScsnco6o8XnHKh/nusozI/KG3x/QM/6wWwXK380IYovEBTLl9po
AEASlnRr9NLjASbse0WTJwKVx5Y4M/XFQ8J+/1cCyDwO7Pd8WvB9qhCbSha4tZHrFqm7q1a7kMr3
NeREouUrCuO+rQI9qWgJhYXG7FkmV6hdYZCRQmSz0tzanbWQUU+0q0EGvJOcY4j8nSCVeHcX771q
zr9BFB2KEALc8ynzbEaiVOsEaWZjLsJokD4fPRYyiDBEIyGpMZBseqNvT3F/2kbpusJEp8zUjGI0
N/b3NGdINqmfCMV87MKOksKAr2f532p62H+5fZDIsabrgN1UkNBnf6cmtbq3FiiGmA9KTjXsYyeh
YOhqqxOGWsLCVHsIMFicTCarn0ntbL9HCpYfnRP6f09+qYcsqyYLiRvtWsLJY9x0ORXXqTHnFnye
EE51+oEz0RzdRLPYFEnPp6ZNupVH7+IniUrOuuyCHlOLWdj3ewQqiZPYK5YeDgkAnKxTmILv+0L+
DQ+PKpF+wIU3Hj4C+82Vld28ye2DtVbg3TMeRCovG3Bs2e2Oq3FIWRq8DkCAEs5mxcUUqtVvbrji
4zlVrV6HC3m6+Xkyk6ZOyR41xW3NuHKgOv5iVgdHXolQ1RLksPxme7vV6pJe9++lirssRtDRDfAH
ijorT9P38sw8wtBBy4aXJWSW7amIFSHJ7LuxW2pZEW/C+AZTmYV+isslXQ4e1TaJ9NGvGxLzm/db
AtRlzR88s5OlHIn/tXDowcS122bfyUitufTZHNJMAavtGfyjA7a4hSgXvXLjHmjzu3p9OILnaj/S
ic10ohDvz+Oczhp7AvoScM9Tik/ql/CPwy2fkDsgTzfSM8yfujZKzXYsWUvZT92lH8IYUbyMpjjP
6p1SRXnSvUZJm372NcuVxGD/WhYyOJHlu636zeDKFYve1/pVwGys3ks2Zm1lvwSe8qU/wjBn/q3/
lMgYzFeGE1zMk487seU/iitqRmET/tOue0TVeOnVyKOx/euhvarLNr+oIiRq2bsRFNOw4XKaarsD
u8FbExFonSOiJgZy5hjZCkrjmynQ0ZJElp8YVHwbraf/WVdO4f9skFFAMjXvl+wgTfPDLU8nUfL0
QA3nvlOuSiKi4lhzsiK6He/eWk2DtXu8Ya8hjJtMJjb7jgCVdRNmAObnq+2CNJ8r9ILKVWRLPLSK
5OsIyrgSc8LrmOtcLftFVAQzn75PA7babx4ncDknO/SzXz5aFo8WQVlYkgmE8kkxHAFAqRCX8DL+
67boiqsRjFLVvMad7srJJLCVXL0mp3FYrAJSbvAhNT32bUR3iXoleqgULrzJasURp5rDrNRpNNW3
e81prZiw9TGh5kloAv6qHihLCqogkjWgoFssLS/xSV4PbdBgPyvuWTAT7b1hNccW4cR//KhQIuF5
r329V0dAIM1KbXLXlSSRBXXzZWtEftbBPq0mFqhQAAhs7GQFbTTA2exuhZRb7bKbSy8cAYzDZQ1U
bIFmq5EOOsTbc0mUedPNzOz+MkihKF4enCNJhouUq4ExaqLDocPgSSxQOYX/z0sQn/Hf767bfg15
uSBj1BKsUaxMnw51jgK04uUxdz8iaZkqv3tdFqtfUdN8g6i6gKtXjSarrTyHg9xkWyrvGpK9Q4/C
9RR+V1SzglhNTXZOMSuQ8PZDeYAYWcDa95tesotDa2PCh8vO7LFsM2J8l7Pd8THLyE407hHWwE5m
P94GOtwDdp6bSwt9T2i0HvGOWP9Torw5NgCCZyg/El7jn7LstSgkpmvJ6E4gn78JX2ZQ4BEFAUqn
BmuHf0i+5TBi8gdN07FWMttoXjxNArc7pgRrDtkOoPK/1+GMoPhPv13hwBoZDUu2O00RG3c+PiEw
p1HJZmr9CnYI0TEI0Go+ih9Tjcnrdrm/rCWknueT+Gl4ci3Q43VRt60kpmFCHwaDicjSkDTKdY1D
FOPAi/T6tbeukGOPFx1tyPnXySVTdeDoVBfkOMquRG2X2SdCSoU5iTWIqjpIWonz4P715jKNpBND
sKLInUkpc5LUImyiTNY9tpzQ5sRnMGRXMmse1XHYvX3EveF1G80yLIqhY6JpClGn6tvrrQcCK3mA
XmjjOEV8nrmkYprQVzzJXhGAKtIHHipI9haOZvBazBlia+TRdDhdPg5tv9Wc62X2SgNXhF49M6Fo
9O5hWRx2SCk5VCD2p9Hz2ksBh9LVaAAqLEqqcyY8uP02e8bbTsjwkDDzpIrUzxjkNX7Bmw7aEE7T
pGy5UpTE/KDby/1+or2JlLBU2F/+vK0qK7Ay0xWCJpLF0kMKJ3MqkkV/ZX2SGMjhEA6nGXusvlHE
i8+YW0ynetSnto5IAnP73lBiyA9PH9CX8F5spfgdpNunS72LSR9tl2ph3QCREJYpxZz0aftxlQxn
PKI5E3tt0jrnnj0Kw+ML41P++GQfWGIGMPaM1FnzFfGcJ7CeUyKNBXjry4eE06/8d6IXLUSARLue
/fiXX0W0IulIhbnY56HTNJR+XHoo3HnKNyVWPNs1rR05gUtqVVRbU13awCXulmBDC0reZHNhBoFN
A7VTSpsDHB4I9+xZtxec5X+aLpriXfUv7IwQYmdS3eI1rtGv64Q/mbPv/XJ6b1LTIBQnkdW2W51i
wZGl1k5MqLJeHOjxbZQ8TVaCwUNHwRCBR7fhCfkP5USB2i1aIJBYTfUsH8Sjn7+1aUTfCxCRoRff
uE07fMHbsJtG+2u25ytCGOTceW2Rmqs7zNyuX3UvppvyhyfSsm8aJCZDHRmWJ+orTkW3bTr2CrAs
g1fiawp5Rg7/KIwMLgZ3oZ/YMh9NgQjx8v9xQ+ewtiqWyT5U+SK+OsDhaCIbW87cYp3jugPJeNRA
WQ4AYe2+nPdYcQMQX2TReX5ZbE8WJblnolOKZFvDeyi9fvh7cnUmp7iljlGK6Qt3zZ5JgpNsx9nR
+yTSKwWpIePdfZgc0tiqO7Z7IfH8WDMa8Ie3dF+JLcmrNUBNQnXSdAxpDw0R+XLSV7ccfJo5cTpH
E8P8+kE5L/029iVFJpRlR2MzYBMjd1VrTH8uFC5V51Fx/jILKJA2GyDTIhiIUEVWGD8eYOF8bedV
QoJq90HDV733E+p42Rg21BnKW+HlOvIlkcHtxozCVEymVMHJ6E+aS1xkHBBShS0sNhT7Pz32+j1k
JxiC23E0MFKR5nvuX5hDdNdOcyUdX7p/Kjd5FjiXqHgucs8xttzXP0jydPo2ODcMqtKOaKDA9gO2
Bh8NhoMKnoFdl7fXva2qqKqwoI7mQ10EFdBQNRaExIV/z3VBPJU6VbG6HH5yTMsHB7UmlbuaQC8h
o1r0ffLAskwOeY0mQ3E8G0WSy/dYM8GHzi5+Li/odPaMFrW54UWvxCNRIYE0nzGFTjYDQSc6B3Hz
0pckUSO0jhS+OTvEcqTFRk9ihzyOVlWdB4G6A0KvCcP7sYwRQ4/CRYHuI858uEfocIok4t9NT0lJ
Ripm0koQEt412Pv07Ncya+dB4Fvt2O/LyENUUU1QSvOBvZsGHyexkqmP8Vg4TAlbta3vN9lDupva
9eKqfMtuqcBYbePckImGj0MKTgBl1Nzl0ncUepmlo/+PYoY9h4qCjvpZHd6SLTgNM7zgEweaCqX8
hsyrzzjy2HYwRzQV4NXknSZnzRbzCZapWHiuR78B5R3Vf0MN5iY9u5Q2hl9W5/yKskLLr6W8wd8B
S5Guha5KWKmT9SXyesC5JGqugWQajgoi60/iOp45cCaWfsKr5IYxrDVQYF0MadRVmuP6z0mju2Hb
g4ojQ38vhZEOnXfnhHkVjYViIUSGp0nGp4bKB8Oyd1z6i7JvC/Irizpb56ggJzjQZH9NyUd4u1Wj
qhN1XGPqamKcnHRO/ZheI+vtTLAjp9VJ/Cm4K+CK63DgdZUmEyAiOgiyALBxUcL/UNU/QqAO+kkK
lID9DprK/Z5vGBu1Zcq0tls7dJVs+GzdSUQBtiW91LJYAY/6zu+INPNugD07X0gRxBJswrAkkLT6
mN0mR2fIO+Aqk3SGsTp0iqVAsfZpGjfPGmU0jlGaQCWjRWqSAw/xzOqTOkWM4ZDRt20RdtwDOcKD
RJuLaYEREgD4+GDOaCxPvqDWB2c7eU+0zzRqb8VLXyhsursb2R84D9w+WmrpmkoGybT0ILuzcpYq
tS3nQRPwJfgIzEd/OfYaVopwWVn2SgRoclv/7pYwPXa0KcXpcNjeu0hGlgu0+C7hfWDjzm8Y6vun
OcMlubw8p3QQmlrLqpCdlrW3LHhO8FaTmms5CehRgf8570TGRcjycIltXc2bltqv4rHS2yYDM6t9
mY61bYFFQyHBV8rYq5C+LevDdxFnE9CD+j/7AzoLlsengKbc8tJl1apNFkPA78NZx2gsfSzBWu0M
C8z6Ql5bVz6/zaUADhsiFVOUQmswwCIndRx507lzMxq+e/eYn+XtIp4GoOruOpLA/eUgnqkbLyql
YzNV1MLRA+OBmk6c8Wu86687quztG/mVP4LGCAIaYT520t7X6zxlcoFv8NC/uuGYMU2hCjSykRgd
M0/DjT8jKBx12MR1BnhqcsZPDqIkXrAjmPWVFUMyUhPWCrzXWXTDLeof/9VjBkJaaHjDz6RpM9AV
uXysmH94zoN3YEdk5LFMdkt4VkAG+8FgbDNPqEQRZtBeOXPdNEnp17VTMVDwLQLbSDIdtr5b8m0M
ArLMxdMZCcgZFjfr9uZW1HV4OZbQt8iZoZeNyf3wZN1opK5eEVY6VivJsm/OEboJ0OFLzJN8in4n
xzYF7+y0bhH3ukypTvbQXyRaXSh+EctkOXP6gVcMGYGDwp/TKZuP52MZLcDZmHxswF/7vu+yU8NB
GesLWbTEmWWfbZVoADDQzG37f4/KInTlEyTlKd63bbetJeICIWKeRm4rP+VJdPesvEryX2L071BI
R380cmRgDs4b5f6Y8VpYQDjEbrR074HZ8aj1LiMSYTXqJDCUWz+ic2ETNEV3wb3vFS3T/t23BaJb
V0kYMBxplTlHejBQsUYMy0TjUaXxkvyc+4WJU+pDSzZK0KjV9RHatC19gFeSwTyy0dlCJnnY3c/B
GWZyJVCDynH7KykwLkJ0/IMel3d5gJKAhAxUHaB5HIrytustzY6uK8OJiVCWCovPQtmuSV1jpYBW
KE5kU3pW1KmHOd/2dPE7Qqbs6u9X8chX4rO4hBvhmP2F2RE1y7LbJuErrXb0at6W7H43tXU3u6Rr
Z0y0vXSS7kJt9VUzrxtpKpryqwfxx/S/7j/chD/n24GN00QCv0px5wTKnqaecDDDOzTNXPAqSlyg
LvOhX9sm5QEy7NyVOHKTVJQT/s8NdvsjXlbizoLCGIVd+yp2L8LD10sw0jQuClnc/83PsEgUrU8D
3tTu2a70pjAfFptE1jJuRiXlPdnNZqI/cTInSxDybH7Z42fC0f04U4OCmcmVkXSrXPobD1fUIU95
2J9wMuKYwbWIvuU9j6th+YqopsAEW22rmLtQXycV2+UzXL8Z7UJOZw7+fJivhpkarklVi5JWsW6l
Ap52GT7+Z7+ujk0kDfn+5i2tIYJSBbq6NnNH8lGEzUVzAheEphp2NrL4vgoLllRyV+xo4zPEWRh6
CxPE976l92FQR6t2QTzJzncJuW0ICfv1QvaPIiY4QDLmLA3PvTpAEkiSzuDK1sVmoHkBJX6wlt5L
Oay70pKoSBVcy2CT6OjpfSSEkz9B3TIYXZLGUCEpWZEASQJM/HUehD1c9DYTPWvqM3deGmlYrNwK
5+nSu7ioYHsAuuTsfVbnu6EDvTobBOE9cNzMslqxPuphdT9H/NoqWCkFR5fnsNbvhg+VS0yrbxtx
fQwyfJm+kivo5YMNCzT8Scs773i/0Wsw0g4nOstk8WFN30rW/+1FOZ8Q+cRFim7zw4i7GOSXf0zX
dQDViGuFskyramtIprPFw+j3MV0ZvRIaK2li/Sta6lbEX69zsQrD9j8Fv7Fw1VGRmVUgFp4QOUID
LclcZFdfkNTtpfGCVe1RpsWBmmSszAb/QDlR+jiGEsOY1qHh8iH0ks6yPfHo14dr+va7eCO3R14q
lJxFKES3hmHR9UEOob7bnJg1Tf3/wlh7KxKM4ai/V0yu/FuOE14PbL0urbEYnHMJH9kytQbIXrov
O/motWLmgJ8ykt76Fj5L58QYjhX1024CFOPtSZQ3n3EU/brxH22tSWka/v5DTitf2WlkAmyaqf9B
oCra4KYPG/4FvgZnlG4ouBigK4ijdSLv9bsMRdxXr2usGfEbE4g/J9aXcMgNyEQNQ/yOywo/hPGs
O1rNc6wIji9ATKhUwKWo23JHim/cTwpS6FKjozmjA7avSLjQdrh10/hAQbNh4Av/hzjJMWksBOZO
rtaO9j+ugAHqAbSeM2AhAbke1XKsM8Yv3dkxnu8XvVvVBA6w0PEh5mLPUXEuh4tFhRGxDBxNSQd4
9lhfzGzJInMhOKcpUWUYEG60bfIfB5/RAj6oUnJXrZc9aYreI1zGYCzLNKQq08gIncIGNxBjnvg0
sbTBLgIcxA3lKVK5AM8ST2+je2dRqvnftc+7TbDljJZPKOQZrquczEeJmT3zeDLDjyuAN2dqT31R
QfcW9nqk8K/kY+bPm66/rOIuQH/dTJ2LrQ+/ABHN0+yhu4U7nTfOtBFE8q/Pno86g6gPDxS143NZ
3hAOOfahwrhjSvqUp+X5Oc50QmZEWjJGeKdKal0jZY3SBR8Dakvxvv3JLaEBEuGstqBpPiG1zWw3
GJJ4xrxOTMQ8LCAS78EQI5P9bIxAdrWTEPbX/cbD2idBwF1tigBw3cBkopLIENch+e08Ppr871mr
hl/b03dWQYj8Zt86NCjn+eTQTdRv5TzMR80RHdIETIr+Yt8qCSNgs8G0BCvG1j0GYovmnJ5jmYrU
EJ49EZKDxV8dpDBB+99nfNQGs0p6luTDJbbacxwBuVeauSErTrAbC00NaMZtbck5aMqBc5EfchLd
LC/w+nuuLkD0ycok6DTui0Qa1gaUDumq6WC41L8Cj+whuUzSVl9/SKJhRaxvCyGyOZ1prild3ut3
z4vypZ5ZICZjXHziHTTGDLt76gECpmwTPWCVhwLesilFYkAXi9nnDCxAht+lREMshY3vblzBXfp/
ejlTsQ3RmMz2zKcfBRNpBOiAoGGwo5pd/O1t+9ZMuNJuFv1JDgAqdFFcR/nMdOX5vZeaO41DWMrP
GfPVf+o1evtsecFppoTwnqFgYWkPnIWBHjw9J2NJKaVRaPfzF4rStJ7qg0Yp0YHiXs0+H9MS0m+l
Pbl57WLE17zNUHSJW4DrUsKI+Weo5kj9VwSO1RBq37988C/RZUOrlAGEM9VhNpofUXbg2HnSsRqv
NAFjAH2pWXGvGgIKeaMxEBkK49bYhprQho2oXpZQK/ZjfTUItXh9Fqar23CfU+9F95I9J20B8zGf
mQxBlk+aHl4leOheioSj4b12OeAHQhMoTBgGOx8at7bF2xEI6Rmd7ZW2O6t7RNrS8JsZzXlsAAtl
CeBLr2CH3PYeUByvWWSkdidarxlu/hlJpD94hi8pqCP6wRWbYCY0BxWl/HwUQ3LixthvQ0Er3dqL
dW8S1r3TfeWTvCKuzaIXcK7FnNOnWlWRDwwcndE1Yw6p3c8whix6/UQ7Hj2lwxkqlzSiARARgMHK
948bYRcj6747M+jjYnbmgjNkuC4V26mBRsl2rwYLz2KWFnxQg31O3RM74ZoXaPLtF/LgViCJG28m
30WrvnC5RDmIR4sK9Sx8dF42GOatBOs9kB//J4jOJy9TDIWdHMRTNTcS6+siZlHbbD0i7MAxq8Gf
GpKpWOLZM2+UOInCf769dYyrVpy8uFsEYDNxBRPVFFFZQdiuNh4xvqN3wxR6Hg35tHo99fSu8k/T
by6PIsdo0yWs4kJycZWdMYhzZmV8engFoM+Vl9GW6oxXm43GMuBNXjGNcGu4H8yBzj/n2Z77uury
YlTTwQBPgvtPdBjhW47bPQhgkFehIdEV/IGpIA0DdkM1LaOLCI9JcxkuxFmfjqI/+bIJq944a1Bj
+hq8yKQsh93X2sF9W9DCATMK72uFnggN/3RD/oFMPv/MD0bBs//6USEVmIPhWHKkH3UYmwdk2e+4
nSvEMew21G2aNelvXcFmOhcObvtKOZD9xIZz3y9v13kJVkY1655jTBx+2Wp7HpA0MBxNXCS7PHDa
DolR3tQu4Rn80x6JUYxe8udECUkLPZwX7OhaZz1AYVACX1s7HfOgesHRv+FWAQWmHCpui8jS7P2w
OLgZLk7IF/UjC5kksH/ceHfIpMVILv0igKoA9nWXQsOxfCkr53WkonlXab2Cpy0hqxcxxWQxgkx4
mXOo+m8/Pr4dO9qWPR22N1nob7Ef6oDyql8lVK9KxbYBXz/e0Im0n7VohoWjN/6V/kMvY3Xxj5XI
++A9dl9F07SB8arM4boefMJde85h2pZ6eBLWekbo4TFLJQGSw2ALQJ7GQvRmRa+t6m1QvcepjkOO
KXrDnB32dnPwjwZpuS38vQNG4oOxiQ0SAUtR/QJ2h5Kxlfqes5G+1fIYsb301e7L1tsRZMthOBoI
00PhyZ+XSS88R+pSbJa83SDLdOMkYS8u4o4oVLGb+YBzSLhX/+Cqo90QmBiXmmQ6Yh89oadQrgzA
hM8g/sP8zz7RvCks7c1g+0H9WB++8I2P67ux00qswHGVkFT3u1IkplZ9gblJY1eVR94URSi1Z6LH
LSOycZG8gE1Xzit1VM6XIIcqt3xzGLpOraaXqNQAR5tAKefgngqzTV7JDjKhgOxjTJbpNyYwdaEo
KiO9z2Uq1nX6As38n1XbXk9hRVram+cZUkfqErOmRAQCTJmKevOYLXSvDLEbGe80zFL7tJgCknWz
NnwcaQBBjYlapSsxqqPCtK9UZ7jQMHZ/of34ArEDnS8/i0fypB0+husMG/HjhyfrgOqm2sP+7P8O
VwXt+/qU4Cl9GJy+1k17E4P5rpgztMDh4qqi5ZXCZzxlpymnNwqPYvSybUD6v2WyCtBxKplWg1/i
vJ/eJDjteh0pTcfjZEjuBZ439QrTJ/amdfCgKmwKJ9Hi+/wqsRZRZdcrkubiYBM+USqHt3Hu1T9w
cqZijJEEA6Z8Hkj7doIeQrr20ob+L8HXoY/4nkNth7+ktzKXRp22VPS/ohdJH/bUsSmoKcA+NYKl
lcbOP7kcpyfcv9heKUYG7+J/5dNAql/T2HukkaMy09KBFD6n75tEWvJAXKFh1os3/MPzgMJT2uoA
n1Q4biklMvJFOlHF4tRmAGYCAYjf0wxp6EjWJQ77rlxzBv4l03OiELZCduMIy6xKYBI8vUiE4Dqx
//Y2wIeM9t6I4EW/9CCWS6dQMOLOYlsPStZpMKplq9JlokgBLnK9LdEE6YcpLqdg5lPorrZKGVC4
fJZJGrFO7XyLNfc4ZyDt9VPyvcvWB7l5JAxOpjejAJNs43yn3ZeLPxnt6Ep/lfNpxudg1M2IqJkV
SGbms3g14nbfUNPbPgkONtFs59LqzXNB9wzo7ezIjDCTmlqwzZGg+VYHxiegkwaKS9dd8jmSE/6I
lKfv17hjsDy2zZBxvlTyRzuze8CVHPEmxHjw+kUen9MYSD1tnzX9+WCNQ7aqaJT/J3q1HBY2nf3Q
BZOPnXfZuc09P8kg4pAZoHraZPnRH3pf1v8h+/AMLd1+avYZavQ2y4Kvh7cyr/OdrqcB3YPOkrwW
6w06zFNeT6FU8czCum5gYAU8HN/zgNj0ckkfQlZKki1m/LQvZbcIHndIQCJPRKOZ80mtqpshdsfa
ey950sHJODFH32/6abqpEZmpYKzY77GIuCp1SUVwfKj674zYhGcNmWgV+ooG0i1VJZXm90wwuVia
NWpcZCDz5034lBnLWMHuBv7IzWcWzOpqXw8aoULAgvXINcXBY38K9pvewyEMm4mgdMAMZCBP6m6z
nqX3tmJ8Q8vdxZdFSeZQIkbs81o5w34A/hSVvkGCEt8k0g+uQmlBObb2vG3sL3C1KdsBLcqqpoDu
qNfkP33U7loGvcp8OpAxah4MGtHUySVrbhnvCJvhtIOyajj7w6N1gPc3N3NWEMYVUnQKDwXpXYi/
lVqRr3DswRIpXGefaGKpTZLzRS05Zk7UhQ9F2uOFUmQk0thKaXYS5EkDV+FRf/2zBLRUnnuKIzZc
tCM/cpt//mPZprTayUE8asCEYGYApybd1ARdcvSZ9OAhSvlswlTKPVAcnL97zkdzBybrTGx6KyOF
mU/o2IxuJiV7RRQNrBuQG+yrORVq3DsKiTlJ3ij7g0HsfYdoUY/SahXFnQqHwCy4EuKunFUqXnvA
PQIy5qTTrlv4kyqkcY/Raxkqt1T0HmadbLqaFen+ylAkRSriv3EeLQLDkhf2OU60inDvG8Ner31G
VN0WAag6HXwgsTRB5orthYhidzkkXt9GJsvpgOsvcskcM3jeoCXelBnmiW8GpwAURogSCcaMEY1C
6q2ZidR3qwTtsLQoGNidwDVMGaah1KzS8fhSPb8SaOlwvsXI6SEc6KRL+94iBf61F1F9asaTxMRZ
U5pTQ1K7zP1ma3i0aqIkJlGlTEKq8loSU2nDIgY+NuAFrgTdK/4VnuZaQRAvYMjHIqN4ZEooEEtR
Klzn5KrOu55bALCXANLS80bXSsDelK2HEJ5fxXJdM7Hu3BOmpyU4yTQKW26cZrSeCG71/r3saWkW
6savYBWBeJ4m8nRZSPxyMPTWtw9SeAuSJ5mEetH9pMnLUFvG6KRsxzDHsDR5Q69La8LCUMqwApd9
QXP6Rd1EApLIBpjccG4Mslkpcx0aN64Br+bQVza9DQ+JEjS8SU2VQPApsepDOtt/VRTNOcE6d3DO
LYUNhAd8mlG140wwp4rWwfrHM6LRw106VKqQAYXdUlSmxKhDHZn3Yr3a5YnEqWN/pMtZCmAOgww/
LjSWgs3o6UtigNw8BX3k2eWvoPKKpCiMBzw2GrTlrH74CmQwP2M53bIhtE1BUzk8nZ6HIGSU42LY
lLowDQNyXR/qtO0KAyiUFs31ZGFlQZVjGjhbvnn/DbEPbpn9zviMk1ZvVMyFNmpctdUqIN7bNFNk
6abyIJftTuRvSKSbbFdw8/uOrPxxMq4KtdXYTkOfeqXy7Lh0Z5WSMF4u0IJaXgLs8uCaDuL15hZF
1FR9csZJ+5fCtbNSCTmLpfArV5Lu4kUEv81GwSab158sqVj8j8xbdoeJDM4tw51ttIp+wmQRWRmW
cFfLpJy2ODWnjyd128WzEbwyTbuyJ6gRk7PvyRgQVhTtxZhQKVgdd2W3H1U5aHTlFJx2hBcw0f8F
hp7q/ZJIYRTy7071le4dzVk4UpcGNsV07B9HiaOBMblLuMG0Q9AYZcdhXB/aYYrmw1PVlKEiKbWt
gAkgKEr9Wci8DNCvT6wxtPKdFNNkl03tud75NAVe7RcKyKuVgC6pm6yoraC2rKzFKPgoEy4CTxeM
fX/g4WnkkFQxjpTNlCh6P9luArBGH0ImXvkve76+JBQr+9f1ciBuSlDednyuFmXU3hTP5I3aDS2a
k7pUWulabLa+OQSz0gQHSzu375aXnM8beOELE97LCzJY2AWw22g0bpbVN2LvBjsyBGprKv7do9Pg
VWhZNajcUYqnYg1TGtcfHwLy3qO6lmAAj0R0Ez3nlEmBB554l69J+BY8oZOveB++Zb8OS/Km5YWS
cV3fNIiRsTflllLHsXUViza2e0zS9CiVikuv6Ijxy+kdI4/ujw/f+iSDNoSeseuy0EG6rw7bUDMX
f4s+Z5QfuCQQJTp29KNCGE0qfmOV46ajDkb3MzS0DaeCX8bBI7LS2eRs2oBEHRYrakD1qA+gnOOj
UZ9H16B14/y+5CPEGL79SJRoGoF4j8oduTfDlQytoXyFAbisMr+XDquqoEpN5vOi9f1Zfc/C+x1S
ZqCdW4Mlejy3Fm6a0EHuJyXxeylRKqzt9bCdRUkr7vfmVxDq8B1cP9U6erBtwywrXZ3euegk0tiJ
VZOyv3wQlqsR9WhKmYxPNR+C/ycc/zV9mDlv5D8CiMzuaxQrSLKuJ6xCarCkfdY6eE5Ftxz6A2aR
ibSzNkFItQ64IehFw0BjZWkNGEpoRG8cH3eDFTXXHJVMYs5KYQ7oo7yJfoEjz2iGEdr+iuZssCK5
/P91xfT6mcpbieiy56yLpz0SIwfzPbmG2Ivq/NU67ixHixLsBfB/wXwofPckxkim5QYHvaAX0C3n
o6i32R5DKHMJz8OYU8alW14o/FSmvk6wXLMtSqO5Nep153jME4GyY4/EbyWI/vtFfUXPdhEQqNUS
7Nojjt0+FwuwjciCtBVCe/1IIgQEgD5ZBx6/oe68furgggaTJaphb53m1umYGO5ykUGyugW1Pw3v
rTxadJhkDQnuNouwL6U8L/+rJwLubdXoNmkbMRhUcJpvbScz/39PiYLrKPiG+TyRyC23QnefsOFg
eiEA5nLU0m1kr3qqzXnwZ35Q1DC+UInRTYfwza1Egdnf8k3jkbzLs2z1h8tGtrADXWTlaaVZiVrb
UjkXPU2uKNHRQCHoEOVJmKDpKoMbZwuaMDE81X/Hs9F+8mZS+JgkRkC1adaCSqJeyNpzc4483dU3
QZ0/rxxb2TbX6PDTV1fTcJJkAfG7HYkO6WO46sKtR9kbnzhTUVEXtaZyqCB4ZddheHjGvJjcgc5Y
rHTMXvjqRHwy+Cwudj8U5IZFCwdAAOlBX/kIskk6tDGdP56PVscE08B8HuTw6Il+EUgKaNCn8xLd
VHWtZZ00Ld3ATtlLWfAz3P77+mDKPUk/7ADU/5xJxJz30AD7sMkXN0gIUrEfLtuNoz54pa0s6UjR
h3IF8h7tyZfAXPXrQixUhcH7WsCeT6QXxv6VVU9NrbV/1RfOwsh63El6Ipaf3whGZ3qIEoYk4T7k
ajtyN/0NtPnfG2Ty+JgSS9Ersr2bWH3XY3iViHv6flJgvWfijkezR+qHhQpH02gxLZPpt3m3f7VD
X8o5MJnNYZL4DSybWPE2Qghdn+OAIZMySCXt20KEsDMu0sOD3nfxQ89l6dI5yAwDITsFiUCBR21M
BtwkuW9M8d6PXtar+yYwIR2x4gYlyRFZdYAF9JoJRgwrfO6IS38kS/KXKwVW/kcZ7/YbUm702tjm
03TmjG1uwcLdAN/uGeZfyUbkbFGzZSI5RXolnhkVsszdaUFLX+BltEEDauEzu5ZsfJuoWZvB6xGK
JlF7qUBUg0eIzWJDdgiVyFmdaZman1RRjJrR2E+dE1zljDLg03Px6oIviV48suYa6t4BDmwW0qcM
MdXtmmtqaMS8+X/3om3gif+aLfbTowvB23V8775wTho6a3uZ0xNAW1vHAh0tnWprhuP9krGQsVcc
Qou6sKfb6QPnAxTktyzFjnPKxuQQDf4OXCwhNvpBoHZglPNaJU9X2Q76MJPf51mmxrzxR6INPmrO
ltJ1cUFVocEKiABAuA12thHl4nF4A7yjqUcvDtkIRdm74AVJaFKM39STPlfdRyvrWUFIJG4873BF
tb1LDwtT6PomAEXVO+dxoYMEn2klRD+UpW7t3g1/npfXF7+KXEgNnJNIzrX5TPTjSS1mMXkr7DBz
Sfwd1R8otp6Bum0c5tITHyM9Zc3jMjmlAiBMkPWupgwSup4G6BrMmZ+rpTXg/mIKLIQ3RAMQv0Ny
Fm5IoTSILZJCRUyh5xhAdfEy9kin0bfU4OGy5Lv7Fr/NlKJhIuenYnqVhA+1ILHaVeEjfQyK/r8Y
sb0uPSimgOvVOQKGqoMWgbBY+98bH7J5/OEStSer2ijuKC928+6irUE43ngBOEQoBNhEV4xdoTqy
P56t9N+WBhn9pQPut/mldYLOyJWSKyk7nNwfg1gk/Ub6fx7sB2oPy7O4pPLDwSfrzikGFdCN/kSu
gSzqf/Q2qbVGh3uDr/h8TDeBJl7whINtGxCjCpeEpQI3HjE72MWHhTo9R3/xCoXoajI6PQrClixV
XQvVmb75P869fzFMvdbWvlxkD7i2Fl2ZYe0la9xLNWvVx3ZgUREMUxmudNE6kBi1gtoVjLHIU60u
/LEqmHbRpxTON6SW6eLPjKNZsSKxebss3IcE7yD2Eoqpnsc+kxKfx8erEIQJfKmwwf5F2qBs89nz
i4A9sxXfyErc7rJQJqVlnVsAEnElm2Cr0gAWPOs4MsuLaAgskmGiHRTQbGfO9UEafJZgOp7PgzVw
Qa8FWaZA8VvC243akSvmg7N0stgN5HiByUCBa+JN5+OOQB/f+Kh5O7yUmCCulGy6q05NTyh+LNRs
fKDuDQc72t8Nr9VGDUzUlKPV9pKHM0IugI96NqMHf0P2NHkXVkcvSJJIkPF629sKN0rCfpfGlz27
8YrfH9spKAbqg+K/N3v6UR60w5cc4bonXwzAWpICv23AYe+jxdKG0CxmZpurlmmDiQlL61iUlDOt
P18G6U8VBYgXTMQzh3HqC0cjVlZWpSlsVfs5L3n8agJICGgk9aXX6SBmRfVkHYpN20kjohTnNXks
vZ44hQlhGQa7fVQUWfDTEYe+5W7N4SvkZlTOX1fFh+xcZqtTOQBpT21QIxSSnlOUhhbgX4EDeU47
jYFcl4WPsEuXvAW8w45XnLZNkPWF3E1RiVAWj/fqc1ib5czeMJsKkRwRk9Vm/PaLMtROktgGhdyk
tqZ7TmSGRZtzz386KFKc3Uny9tiV9I8aZOlpGSYLExDEGjvU4l0E0JrMWFvTDrL1GAvZLlr/Dv8h
rMHRIfbqQY0M/JbOIEbRCBsu8zBsMBln0zSeKn1bufyoj5fHF3hdkBQc4uRP8B/8YB/gNf2cItR+
xKvSIWdRMveCaUfD8HJT4duOKlGAia3BJL8XhG8Dn+s2RDakC3PTUrlWRHTWGR881YwsGgtxtYV/
Del2WVSMAyGwn4FDCXkIRscW2cNFKxXy5JZnM+K3OSHPGDv3BD1lc90jerWc3cgoHxYKZdVmx5nG
Pk5U9xPA0rDEKFwluiO5bls/X76LrWUY699R360MO7/g0qhC5UdcGNytSWPIZ7G0UtQae7Db3vJC
d/swSg10C/67t4cN28Wv0ktZSEOMayMRS6/1UlwoB+6JFi+lIQZ1VxXyrq39jocaNMrcXz/etXUs
htefK/Bn+G+2Uh1psY3N1XGl99QmbYC+szeYC6MIySwcfVf9qzPV+ASDkGT/KFwy4Ss2F7Ur+8rQ
4ygN3Z7K7+XIaKL7jAmPo9YZfcxHz6rGWuLbCzgA4I3EfYneMLr/u55EVqWRtgrAzty+IQAdw5yJ
ViUyposf5ml8jiq27wTPFGMcpQrhPQ+vD52TqaoMerxkDl85+JDXRYuzpk1ljkVm8E/kO3eGShWB
N+7+bIGopJxO14RiFDJDFwLf+x5h02SU2167UEkmn/sn9+ntutYPnoX4mLmjK2v/ONAqUcmTvUFG
zzJS0nlBgnMuLEzc+yzy4EARf9YW98p9S9lS83nYp+F8IRxXamPOMR9IgIcCH1lomk+I81jUKA0h
7v8RqZX8MS4TqH/FGir76nzv1dgJ6RNeRNyRtimnt7gTUF1BDQcxU1xTNwvNLLZch34Qc9+gAnJ/
6L1U7cUE7BE/HE0jsf8VnXYYVcL7nINcIPEmftnh/ViCS3YHwcE1XE+AitjDXy1bKFEMJAwimfkv
4iUOt9jlbUhRYx2N+8IG7L+bAr+S609wrCzFDV9P40RZK1+UAzVxr/Wv+68EBqgIqwytBsIEv5bO
ZmUeX6MO+HCV1cYpVpOcvbprpl4Pzuve2L66GOWQ6tC36pjUnovNC6juWxhkKeodtUFd+DLBKkPF
F4CXvccOhEHUeBaK7IX00NBffyw98CGcCH3x3uzmSxhTF/JTToQZIq2VvBXRDHpkVBGeopMR4x5x
VzMoxftMziR3U21v8fInK1LPi3ZWrxyLqnV4Frm+eVNCl09xB1pLmh1Fr42ik0sOuku54rkfGKD4
J8ap68MBrP6/B2hx4W9L/QNe5jr37vox3plR5lLRAtA/XIL63945Ddtj4KyBPLNpPMv6RDL3uVoi
W6B2eoT5JsBZHzrOoZLUZiYTBr/tAoEazDCsj80197xVBILHo+ym/mRE2o6zlQEATHd8GJQWd2pP
i2CdK7yLGx6d2Rhb6araR2Tx2PoJXTc9F006djC8r+qYwQd13ZQ0naiF2cIvGY72BL+xYJp3huDy
5kegh0jAsYXvgUwQNjA7S4Is7RByTHqzKMmxLG+UWTiO1CT4lXWijE0HbAYnYb9JFaEfbK5aXI9d
2IAG7F9Yf/nWt1kd1lQEtfMniiuvIHHPm+S6ICfyDhY+GSWY9m3cUYF5sZdvPeO8NnvUGbBlypY5
OssiZcBPn28Io8hykzPzrfmmMK0A0Kr0uPooNVf6+99491iMJrvs58cAkzHMOAlXKrAseG7dFUoB
uSD0cP3RmVOlOnVgYGzbDVxhV0wySBgjhgqSGBBnMKS+bhrCAbqIgmi3GB8+CqvNn+4C0xOW2RE7
HIrgaz+OCeFemWVHNcj+XWC2x4ySKohaH/KR9n81eafaMD4nEbjnDuo3LJ6tE3DulisM/E3+a9A4
0HBTguajBJS0qCJmRA+P32qqA9HO6R+5x54ItKz1LViYVp2aJqgs4PJAx+nCkpxfS3fpEC7RsgfK
qVb5Qs+Oh0dpcCLI567FjfPnxPRFGxXODs4v1v7S0CGOwOCmhPv3Xqi7BnyrMonlENw0jbUBbk0p
XXbgXjmqH6Qmmvv/yr+dk4jLL5KuWGUfGXZbCwtEklJSQsfWXkN6ieLdunAnmgbec9nWKRUR1Z9S
bj0SkPwIFIIzcNMNkKF781a8AGfZ/Xbj9jTebsR48ArM4w9Gh0HSFVqq8+k3KmKinDxKgCm8gFyF
mHEfrgeEi3Bk8n18s6KEvw4ixYB49FG5XQut4VvUlkgM/ieFZ2YdASI42T75P7pw3ij5L3y0SWxa
XAVHq2/Lpy5W0mEpNTyKLnwWpVr88j7t+Wbd0bpZS1ihFUIi4CCCuSU8EOskgtN4pbdafrDrfW/S
WuhxQ/IJvERfC7kan1Z09OWgoDY7Q9n029bz0GmFSoyH9YXwLff1m+mxJXvXLxJYyytKr6dOQcMk
az8JibAgTwT1wBcBYnTPx0bImwEt7CvdmHr0thDjGsDchbHkwDopXDPRDfs9Pnn/vidtpe8iJCLg
FwHPw76WKrtPIymlF1g4D2M+GiaGSWDvBFzuYySNA1QNa/AcJyfWCGraigKdJE9fVZ51312jgMqC
jm9cQ/b/A05detouwhcS4LOhxLESMVije7IAQQZK6QnUiQqmcyB+ZMxwaHPnTgc638SD4nHo7cSq
mDvRa/Qu5AFky6KPe+hle6++xOSZmVTPH8ZuDpk94nU5p8+d537OCnzN7P3mcGeZ6Ickhacwoz+H
wtrgPPC4fP+REyXeKcn613+jNWO8yceB0I0VtdTcTECTUXtmkxTE8HdJoLg16iQDdk6iAw2Ixyl4
FLPYlW6BKhLReRIvGWwUTwIKBgx/oyUDfelCsMR8kgC/AB8K3gqvUr0vqgVDc7Qdxg3UsLvY5Jzg
iPqweCW6tQTr4i6y7YaBsWvA71omQKZYUrmT+hvSEbo516WBBeGi1sUOVdhbAGbWzeBpqxbt6XQD
XFChkCwrGjcFF5ag6J+5j1jG63+VOqV0tk8gOOSVf/AIx93qTCZpwv8PovSzLRBlvwy/RclXNYCI
B/taCvFx+UZ33l+nhnhi96Dmg1NR8pcsq3iUCth0lB8/tKgdXSpC1MBMdBAfp+XWl0QJDoSyLffs
m9QyGSbxDbYBb1hUH05moCG2sQiHxvd610jB2IwyTapvkJX6UNm5yFoc+eLC7I2APxyk9WfyOEuP
OjgJoetrCJk9VJw+ciBaUSVnvqW4oScTUi1qnZUl1mncwYwVf96SkoLmwmclYKgCKS71CjoBCvT/
k6YjK40kOwGhKl/irx0MeuW78hkB6LdCbyvCeqXylmlUFkqR/OUmCDiiT7tInHIii6xNj6zU1rHm
SN+xxA7gncUpugQvbHJWGPlIo5rdAebjeyy5+SATkYKVDkN4yWbMo1LxjjFBFXD2HqLh3+9O1Gwz
OEQeysmGNsJtqbATPaeXcSdrlMmeZ5FWYOi2LAPf7gqDhaY/OVVWAgugrr/2vCwtHfqV9S1RgcxJ
T1OmN8ugqJX62xw9Lz/MfYwkR4G1nDr41gcJBMyHaz8PmHvRCLm8QiCO27gXAS0fb8Py90LZCc5e
M1ODC8HIi3a/0izGyh33iKV+/dtz7Rq9A7dmLNAQh4fam+6kpoZ7bDeCG4MRnuE6ZuOIglEYYR/Y
D4OUo+yFkOWAO8+0oWlgQP3GLcTnTQCN6ucZGy3TBbwG+9PbUJX2yvQ6j11eAOtCokYZogT/YY4F
uPsoKS1n+jxPyjkyh8Li3QnOIVeCcDCNwO2OW4AE4iugPDOqSK1wJbHTS+5Ybd0iKXWDZ8m3ntEw
GqcKnpF25CZypJaSvxsWbPbFqJXcXDoZhNKKcOoIi1UCk9qpN0XnbsBHNGCUeX1MbwNLarPnJktR
sV2/ptUsN94XBHkTO0cf9XYeE+ANVXcC0i436UvYpU61rTWnYyLxINnrP4Ejw36bz0h4n22IkV6J
7z1DyMHuSt1is9XezKhiO/0d/YNe0XbhW0todG27YYFFXL8DjeUCV55SEkExJtlwHbe9z0njY1ju
9UlALLMrYX14ovHJSb0FRdG/RHdkaM15jIXToTWnv6OpAQmwoT8YWJyo+POAxBgYv3xDlHc395LD
pvn2UtTfDXp/69Mh1U/Uq7Yb629aBVJmXfWFrkKoxFHzGMwrUjj9Nlt1yW6eDiYxA8kZOjcQ1LBO
/2VbpFiwSpsZunOT2zK+NjmChQ8kqH7mQhJ7K48l52HYuYLxm8XFSepO1j34I4IHKlad1Ux4/JmI
j0aEzsahksGcvlKs8bkRwrORQDzY6PfLGpodmL20Our8B+Sx2HdH5ZoW+ukyjigFjFg4npcA7rzJ
Pwme/X8wMYsI1L9gGhrGnTTVS8KXbywz7XUoKhXijaecbxSkBAOiE31H/sXC5tkEQwYuKFgiPifL
vIV/QVi1rvyG/PsO/mCqfU8sMePTXG/8wqHrGQIlDDTpueWnht7kjXFkGqZ1fuNuAH60tGe59LCp
a0DLAdlLfAfuPTirIAjeOt+kssQdb811vg0Iui4o1jjxTUxqRKyDZuHkPKhWQQV5TYcILXRF5eRf
xa7jXaqMIyq21dJ6ig81aHrkVuHOzHt7hWVCF2R17Kx+alM+IRvDwwhET/paz7QB+S3Rhm/6MTxY
GXYF6Ehk6VHSMajqFzk7TJkRwLO5PLwRybkEEvailTZ1CYZ26pLU2KKJ/bgvZ+kt9YSSNFgcjNAC
VgMQc2LrgBr6hbLlKoNMxV6kWu2RRb7B24tZccxQoXS+f27nOZLogFgOENm08+Znsl+w+Hn2K9kH
EY4Fn0vh5KJ96GzEO/Camv2dJPGubc2Q5xQPqUmCfYRaqEnkNHKdszp6KNZgYXl1xdx6NwI749BB
61BCYnReAwtZ7UHKMON34HF5Q38xD9rS0VcWu9eSR4w7v0YUWvQ6d+7V4mG5irnD49gd8e4h33EK
i7VdJEU99AY+A8zoPXIJuhyydTuigc7cneK0UkOoqkBCkUHuetvkk62zZVjEZTKeAke7QaC5e5pb
ZG6iKSi7P4iSHUDkx5n5UvitEZbR1dAezx58dwD6zSfs6OP9/l7TUcXuBBpvbmpRdL2AOUXH4Y0L
za4GExfPeAwG5pVsszNUiQsG/CPNIYPUE1QMp8hxnXAo0fKujqqizY9Hb7vlmdXi2i2bdZuEl/V1
Ui0T0Bl/i6v0FxYyiGJRGdgNxfggSWfSQzKeY38EcifZuTe5zPjskgw3BP5+72SBdINb5e2AsHpi
suVthB31eynFZTNlX8bkXBW4vZtYeAVjcvQPW01NRbqi9+D1eFlcMJH8CumtuW2h2cSkm1UF5jw3
slqHn+ThIzKidupBXuoAqUoGnzvJBwMch0SEMLIMWqWxAD0Mjlo14ZoBQIbmylZIDy+r7efstCr3
3Gmymy6XAjNxBntu9d3A/F94HHgBgq5OvQxqA83DHAhjsRIDbgyhIOScRvAm4+IVJPLMw0vZ2ycG
S+0nP63oaQyCD/LvIfy15/sHNCBX9ku+0CjMl1lxxpw1drDjN59v/v6Hkgu6M9eDCBZ5TEEth71X
swIGvjzsdn23r6dtpgmRD7JfepfK27w9w+9pL+8S4AOr03MaDrNA4kN/1/IQTZJ3T7xmaYNyYicO
6TkycC0C5ARb+fnNHGeIlEyTR90h87jVKGtxtig70MKzml3bPJpU3UoSVy/FPdWpRFv+koIC5TKE
Xj447nX3/KEGVJE8nAxZj0h5FoB2g69EV8qtrjylZ0DgO2Nc061PTFtZGjWjh5rTAefEXGq0/8of
zq8cqcv6pyidnrQINMg3ldgTKqcDV2h1LnyuK81lvU8uoKobM8L6+XCY2cr4v3cM4xaFl3HgpSiA
wEqe+RhI2LDJlDumJBpjUgthIiNUrucLefMAIPRvrZj6E6qv9CKVEmgT1g/cEZdIycEMlvteXifJ
rV82CT7Xw1bMWadl/t5IHxlsT6qU8Ie1CiW8Rz0gn661XSk5EhvYxZ+EAxlgmzs/gwHI6xUi195Z
vzJDEKExzea9LVrZKceJvJ4KkgMx1mwPxX3Orx+ieJZVOG3+3iQFmC0jn0fZeeLG3FVYKIQ7z6s1
yaObqDmLosc8phy2uUFqpmiao/WoGETbUZHNdTM6XyP9U4a8XDnWksyaW//2LbOWd3v7FsYUUUHT
zeyHebSffBeDDHZQ/KXV6VNpbOBY5g/lNVpRsQjZGr984TX+mZOJb1c4lSCd2du7IePaDtMEhlTJ
5eeGWXfWDK8gh0UdQBjrjUqircDShgpG35FFWNXldXkaO/Wv5ZF5T4U1ddqzrD8YbYhIpqyKwNAj
Qr5iItvh4J1pD07+YrVd46ZRxyPHFvyE5sUt/QVSqQrr7zRpaNmUT7Liyf4x3mq2VPjY1DGFbzsh
6G7UapgaMqglRwZ5NKYsfjHpuiJJCK7O4WJc1pmkwdWk0i4s6tJgr91VfXpowctqqAT9M1QICtqV
7lL4DQ6Xihw3tHofIZyNoyZjknFgnN8SCOgmOkJ7dbF59YKZL7Kdcr5IzPH9U37s0KrJZG5VJB4N
uAMtGPugCy3Hx90Ud6lwRTE3777AXoOzEwqkqY+vKga8jlOefkrtvVqScGdYAt/gKdgK3kDYZ8QM
QrPLlfRxJQZSNqQCdcku7W1MHiQsPpC2YS+M1lsL+M22LjZgkN3upfehbvFnIekTaHFA4SbRnnrd
vCIWeYYZL6/w13iOtxvjlt1jU43Fmx1ZJSYaazk9QjFnG8MFdxBZ94KbrhrC09unVl6dQL9gXjtg
0nYaTqfwCkWxq6NPyGHTcJM6KA/wLBYfS2SgMhO5wY8ykHQOxybrWXyq91Thy0tKA1t0//7PW50I
3+z3QcYlMZxU2HFvF5kV2fROhig1q41Nc82NP6FCgrEbM2qA6+aaYlJbXqMG34gMoNAdCcaa30nR
DGAph7RdduIWp5YTBFydfXMTlGi3bqeQk8ONg8hV7OKwyCeecJKB4ZSkjRT8sQu9ctn2Xzib+e7v
lvXvggTSbBhyinFIsIgm+BKS89yr0NEgc4Kszx9MNHJMkDnOenrbrQJooDrEyTHcptHIUQpQ2qFE
a6g15AvJZYg9+xiUIY8UemIOZiOB3txI6f72862A6UTc8iVTspqB2CNM4jP/tcjeLac4Nrnvg2b7
nzwjNZ/kUidxYLhaqh5kOTy+UOgJ1p4PwBtG4FaxWDI0NMtYQ3Rx97oamA1utIbftGjDF6KX9mnp
t2TknHjRPE7EVqINXyk/00hHCxb/CTFj3eBhOqpF0lVsfqRXZgVNgKEr1VBjoVhaY7Z+wpemLmPN
sGgGCoSLo29q/ZXpmbE9PMCo4jHwQDQe+mW/9c8l1hjtU0sc2ou/kGipqA3E3Ffh6KWkXWJguP0v
b16VOP6GvHhVBUnVHWYYhBxwygfvZvg0r9+H/NfRupshvWaQyPDdDMQC314Xy3gGjIrUXUZI6zTA
vFIGeUAZ8TEz2DbpCcb3uWQW+7mbqEmTEWwLbgz+puXWXx5BqflJlynldpeZbOB45R8Oe6RV+8Hr
Hz4oNbyBt585IDGudjJ7DmgTCojmH0sBhu1CIofPHbOpCrH+OEtp+huyIvtKqV18Acr2AcdPyFsL
cRUQKncR5hv21nvS25i2XDy/pbgHHSW6klwbIk0SOnKX/ADFUGuq6HpfWUaCUIOhFv4mhe+YxWix
4DcLIzSs+86uq9gFZs3NytKQ0+axt9SU/hsEmPjDxIu+EOQpCRUNcEJdjCEBboA5noaRjoA1lbkT
y7EogNUAQui2Uktwc9hmZI7ptSnhrnSq8Wqk4iRpXZcQ1gmzyIIHR8bUmk+29XgdoCnvwBXqOoYF
B4EJABN81DVK3zOe41dDwBJfD5GNa0Z5H1Z1sMLfysQEn6By2QKoz7rNWVV9vyRLp0qaxWUqCGRH
WvhJDnZNF3LxDwyofMblLkbgHhKY8/P3Dgtca0fJnJOhrbi3RYiD0aloLK3XbjrQs3Iy6yVgzHMG
juQtlULHL7nGzOQuA/9OkNsPHQwGEifMkTWtujixt6wBnejaH5TqQtxBxxLmp8h8zKmdpWaQ7boh
W5S4CwBfG+1NatWX+cS2v58p0m81OfnNxhtE+FuXM5rYT0xNBRLr/cBu9Ezu7mYJl5yBfD+ACIuw
9cd6eeetNlEPf3z6ktja+TL61G3/PJrJNp8euftbNu2IhuwrTB6udg5Vm9Cw2o6ZRBDtBJGTzMjy
Mlic8+W5WbKK5jtCWV/d8+tZrMdfceEbYR4aD5yyf9CeS09RybvBQGCTcOKyMoGy2OID28E9ZXu/
ibjgFhf49SLSAZVDxuILJDutoguCA8x9FK4fl3FGO3qJsDYGlpfTpnS26gUGqj3WoyN4/a5zO1rG
46yesrzWrCHhEiu/8/cLW/QjPl3YfHCQW4V4XC3xkPoKE0oiVr3u8UAb5b3AgLftR9RJIguR4mlg
HzbyS0dnhVCvSL0Hv/2MVelVOGfGrmbDIS24+bjmLaINxjqIjQ+Ups0yo7b9YVUDA5RRR+Q4IWw1
1oiGYJiqOsaYGK053hr2g9UvO3d31jQLNFbHrIXasTvJFHa/xipSwN2BM31y/+acVg7Ss6O11NVn
kFdVIDBOuNpmHQrr/jDZas6RJjRbUfyRWwnuDH9NEv6AQut7DluN18QI1ppKm8HjxU/TcuiATdox
8qGRVguG2IRCZvR23qwW/jLACHcxUXq04unFpwTefl01MMr4NOC5tdKxtmTyg07n4n3a0YuMLeta
V8C8vBxPKZblTnqd0pdOylvMk+6iR0Hgzn4+r/XuKBVNcfKZMwJ5CrdxrCo7cjGqjyvyc8CgClND
AERUdc5hOZX/MMLdWML4anz/zePyjaqP1MRRwXienCKQTRNJ7LC9aKWnhPjqq+C1D3heX4zZ6TX7
SHT1bE4tu4gW7WyKtQkW0obu3mCLV31CpqM2UIcJnzvMzD643n3Y/+tu8oUofOWllJSw3CdvxXm3
81RZY0Fofvtz/BuER8qfKoQFw8Pgei6ZIQCcdV/Nw+UYh95epS6p1fIc9vhDy55qQOWjjL2BMbT8
52i5nq0SVOjWLyrCkRzhhuTEuAo3GvYgbLS/vVWigu9V0m2Kc5pQOD668qQ/85dhVY57U2nCML58
t+M8rPa9pjw19Fas5fT/LV917KnXau9TcIsrK71Wl/9khHv63SN+j1/9Bm/w5PAQ8xLAxZJeFUZa
ji4Y6Jcs3HYSrMDGMd+1D+44gtIK0m3vOuqPDbDM3o24vhvpBoDDmbCp02nPmX1AqpLWAkTlUYob
bsjnE5V2wAsGqevdlyhspqr3A/IpY8DFtccwSlRIIlF7F7jMenvRnODGCWhJZKYmHP64w1zWdDzG
je5Cx2nMOTSelLtVcj9Ta9FVwQBXWg8o8JYqLUfDmEaa7NskC7PCe8r6t3sby20rF/g+4B8pmO2B
ElmCBHXQh4XZp2wab8fEpC1Ro8rDKujH+NmC6NFe/cniHLwQTWmuFMXeZyt1N/7G2suFJNNkGTpJ
tAYqxm58ZXyx0mfD8fdImaEoP7AvD6x3DWiAVlR0bVBFtjDZtApQepZwtm6UAvGKkhnmFi0PoFkn
v08M6RVpgHwqlwvK/n2W9PdSO9ib85+Ch4wpbK/6raC/0Ppw/1gkArg2iZBgeaTLegpu4JaWMfZO
ifhfCvXyvpdEkesuWdDn+lLHDF64FYRyQGkiF205VQDDaVZbRO4VI9YOIaysTFbjgjDafKZTGzQz
WhRiCjxQH2LjmUs3+saYzwmGUQZHDHtcZrNxU6LpT/y2Qjlug3mHBsOUkN8iBksamTwkQ6WXfY9E
IQ8uPPr35sxvKSHt3ROnV/tyDxARaSgyd/RDAd9LUzSVAFxO1qvoien46s9Qy9zfLFbUujFsxN7e
O/v8e5xQxpii7wl0d+lHvwtBtJrvtaeWQVV2ghP1ORDn0uPk/23wZw/SDlXYOaFnz2h+Adh4uSr+
3oKMzMCfybXAL7RBHeC48C+duU6iZWg3BrNHxumdVPzZJXw8CbOSn6qik0KngUqaBLTeJkfsJaVs
/GJKfIWxk7vzmnqTtp/x/+MkObnP9oLHYLVmzvj0/clg7lKR1I/GjJ35p7ViiAxam6q1vdlo/CRi
GQe1p/44Eg3mL+fxAPjyciPmdnSJ95DRumkRB5UMkpMywcVyGPtmorH6E9qHo9RGd2IHwgy2tXV9
aj/WtiQx0WD4YOiv+uCRFxiYWl3OtAbzkicI7hBWWoZzslv2zuWgrhccXoA/tWVwZqeiMLCePGu0
PCzD4grR1NgUbPLTIArJz8dwh78dAWpmFKi4nZRJmXw+0GupCz8W1m0czojqVAnqOMN2xBvGJ1/P
ikgVB4XkyPDDr4Zlv++na72jChlyE2QUHIXMCWax7NZfZwm1JB0mZ3vLhKcwm0049xE9FkmpTJKh
15qUfhkr1iMNKJZuiFq3c/nL8o4eXrRbe8GKrMvXPnPWvbSn53QionWvN5Ly/iRh/ok8Zlz5UmQ/
45gXAHfTrhd+0dltgLBYvNOYiDu/+EZOFa6V7FQYXmukHWqyVxNNWOCKwqKs7M34yPvAiHuOd/Ui
BTb1cDAl5VmxyzoyntFFKohGy5f2bp9b3tjFrafLSUhN6tl8FpY2HqtItaYLwTFaTtY31yQIUSDR
7pfZeKJMp1Ho6NBccS45YmQ2xNKoW1rNG9JLolPfp6hedx0RaTiWq7pRYvQC72M2rTPbQlsvwFFM
9cJtprjxe8khqFrJ2aK6eMvLFCwwzl0DxmuCZkmIKgBBPTM7CHiGmx+AP2M5AzQGV2dQUSSBBxS3
b5RKWKjYLhS9vLf1xfu9fGm+x9tYrvaQb7oymKx5BDwHTSRD6CrpOQMwXgiEpy++5tWMQSey/XCS
p9scuya075N2bnlkZfxtykzk7Hkf1INVeDZ+GZRob3JfRglUrJ5R8tuhnq+EWnojOM8dFU3iGIlh
T0b3148buYonh6JwhbS2fvYIJfY7vIcIXKN9M9jVDWrr7otQ+yvREQecfWTToLiPCrJ+r63pU8Zi
AtQ0MSm4pdGq+LO0BKpz8rxhFRJm1P+C8oB9Oa+2JBrowowKJWG5OSUVhqcmCp9k0EJTd9ndRAQ8
lJ464pdngVARrR9oJq3jYxI41mTaY/Lrj9jbKL8pIqFUWsxN2CvDCH8KomPxc6X/L3jhJB+OMeNs
FA+H3LJsmrPQ34kcl5HBmyp2F5JPGswEQ6GtkcQWWVd7ZqadvdMLTnJu9AzbQWk8xpvMDCsmW3q9
XTusyktT6LDIc+bODCjSNROhtdIpBLoSLap1bv3/o5GxvbRQKwWVZk19EVqFbw6G6mMcCEFHqpik
Sq1QvWlj29FEBmb+A5M1bhcZBhEhJ7zwDRZEv6WPmTYLVoKilj6uaivCeeIInoz4RzSxaRkaJ7Ai
ljDEHXrgBVeISIBCTaKNfeb5JbKNSeg9eifW9udfHB6LoGvrJ/d7kCVAQ1i9wity63JOISf9vVig
l3H64KKfn6QDH83HZ7eWkzl6n2sMZERMZlK+ahTpsXc6Ra+4/vsbo1S/zIyPkJfkZ01XygoP0yUa
2wd6GVxaBlE3b2bOp7g4sD92yJnH1ONiCUBPEFQzR8jtK3GngVjPxxQyduql1BhGJL6FNsGuz1I0
y63869Ca3DtDNeJmfw0qaDLtbHv+HwXBhrhS/h8+zuUIKyUy3v2SgyvRupqb3q/yfGp1rXYFNtLL
FJHKphhVFTbWDNfzOJj776XOcov1GRsNSwpdAtzTcOKvswq15e70ns4xvGHh4L72uIRJBsG3R50g
eJ7WGxwNHu9LP3WoNvn4zpLfybTIIOVfqPx6rrKj2GWc3zID3PH/jL6cZhH05FFYNcwgkXbk6TeQ
553WWVpyQzCy8z/FLkZHmoEyyNqAF+vSqK9VFj1rkL/p3Ii7Gt8cshuszXoPxZPnBeEkj5fUzEcR
38JEsL85WK6tMfl87fOY35y0P/3xNHIAMfOImtH9osi013llEUZ/6G3mGitwqYzD732hpBIKmmFb
ZJKZCgXGY4l5ehNzMoeJdJ45kSsF4v2mhXMojrx+Er9th8/SSHz6SAIgCyvV4vYn5nVO4oC9BAjL
ebRFiA4qS+w3BHUPBPrxHcxhplDRblVm8J8++Qx4c7fT6UgTAsCMPZUvHX36+MJQN3L4k6/7LpcL
9mdV9FVadYCTDsi4deZjKMDcVMiGmu0C3O2PbEoFv9fUfsjDC5vjXjs+4Hmgs5LFNqdm5Fo1B+r4
jss+PNQ0aJTHQuNcGSc8dz2y6WUYRHcrxFf7AEleR5aXXIfSCa/+pgqBQ5gcRL+TokeY4AsLMER4
16CvoYwY4AXZ1q++w055IcnSvZlbU6kndkrOYJ/E6u/QXqTbRKFm9M2lc24SuM/JfqOG0ADPhw0N
DqLp+TL2u774Dbw6mcFC4+1xcF2eD10bBwXakTwFKY2cRgvuXk2rowGWinIdoWmX6dKxej6WK3Jt
O0RslfJ+tzgrX9+/nvkZSaC2j1oEtuNvHomz0unxnK/WNfFADt63cSqrOW0PFTwkG+C5ZoUHsTpT
x76zO70EfkHpPdKV00FDz/Ax4glCcVsRJKPIkLjmg/aHVsD/hPqPZ0Fc1KOUZvmVtk7J/J2nC2ea
eEj+ej/vMLRthqCHMkZstdUlJtuFHxWiJTJro6nKxX08SvabMxTabAh8bUgPLs5CNsUrjaY/F34S
dltwjRGitO1v+XigvpqCDGMwilbV4DLluZmdfMSYSFL9M59iapeMllt5MAurKQGyWu0Y/yGpQVtQ
GImlbA+fQEoW6u+wjIQbvFQCi6GurWNOK+9Ze0XMuo4DSmMXdRBjEyHzzHIJ6+vQE9jXyWUK3ArI
L1+GkSWpyc9EoR7PG9ldfu84VVMjkaa6JDKRuEusoSTcIRrgEu3ONhNwB8VkVmln3N5fVxa/xTk5
r96ZR7vWnVtyOxxtpsrLdzK6K2ptbEUK7ewSSPymZ7SX00XrxXmdXxe3xSArUlDTHAlPASZYB3hQ
cMC/93O5lvhKCXaN8vrjoE0qzalGm0GXNBasB3WIXVUWur9Aeg0FjE6KNlPt1cbvpOl55XIzL61g
vIm1VWLcpvpqc83sbVYgU0Ar1QRjPOMuAeGi13hXkddB6HccO0SOge2TPtpIArYy6J4WAH1mcN3+
TgXwPQjnXBRvcs6Dss/3zYpp4yjcSz51pm/A10Xh5Y8naK00pnuRep7nLFyxCHZTOyBHTBri52yd
tMKpV3QNXZHPF/2whMKISuvQ1KOHWZC1H5YfOT5lpQp6IkBcTfTtfd/WpECcI1KgWhpxpVdjqA0I
L2juwApzmrrlgekQiMU8weBLpCowibzpmJ3E6A+pQYFHdXH6Fnn6su4GDhr0wgMDjmH97pAs/Op1
qUh8y7vaOaqPjgy+xlofsnkKCXlyconLHGdBT79vRhHuFWv6X9UrmXW8RDh06SVh+fKrpvRo0OBA
pnUVd2w77D9fP5E9ejLjCOublZGSjYNMiqv9aKG003RWPEig1hxH9rby+EskJU9YHW4TWGTnq1qm
7F3gIp/UbpU70GB6z5zl8wTbBaPqI2k46cqqM9tJR6o2OOLur+OwHeK43oXSX23uLmpBNTRlJ6qh
PEwwFQF0mXkE9auhrpf9g/P5sDEg6k48j/sUbk40XfsgubOF62j0pfZq1kto3spuRnDmrjtFGLig
/AQ0Vuit0uA4VgxORynDharGezxxJuA3pCQ4XzS+68PJ4SjbDvc2YMpOGBnhF/9NJk5dbWAyK/8D
l+JRnxd4eYiwQrK0/qTdf076qTMtvGMooqLRd52w+vdr6F8o0trR5At3i+9c1Gpbjr/7JgMn1ln8
ucbE+FwBql+u7QdAZd+epyyByzm/KqwE+S+p0kxKnJxeAqNcsug/+lez8K+qT28G5cTr9CtZ42Ev
iqhzhfs3Q6orMYJr9MKYyYRAm4cxn6dNSmkZIBMePHBbIrGQgb3COJlVL9f20e2HskeTFh0T328m
VyWKZhjDFo/RpQON1vwN/RcNCN94I+Mf23uy1XlpDyoYT3ZQSVm9erh20YJZSReT0pnaTouk6Xrn
wB0gRiGRKLJ878tMCNUXrnT5dfdF+1SiTZ0bt9oULBgN0ZT5Zr9RdrXRy4lamB0uzlNn5g7NsHx6
NA9gao1yeNZcqcNK/ATVNQ8C5xag1q1OzewAXEoRljawNr8XxROT2UFL+sRrDksXosl8eSQaORfc
J1MDpf5M1YFVscJHsz/WT+zO4CQ8pBkG2y4pc+emaiw/EefGKw8TlbOiobT13VLxKZFrBQA3uomg
vGWyenn0ZfBWv3Wh5ybPW6bFERNJbwUvV9T6K42PB6ensxZpSgkRHSFzEKwUuPtATg/FMXnhX+EA
tLt9VRUbP9ocHUb5hctkFds9QiJIx1Kd14+YLezeRbHPcU0aaPbLPEe/XDzJLERwIE2P5lTAiNNz
PuWRLdgW0Ekle5nWeiH29iuZWy65mGmWm9rfClHbWthcn0EE8z41liavhA4BbxnFAR/5kx4gXSMv
VYNPHmIKEO5ydK4tks4m0L+A1hLtUtOg2Mz7UJZx80BGtRKaipuc2QbtYNejyGU4VrJc5jF233MS
CE8AhxkMD/GYk0/AcRe55cfF2P9ij91n8BQqZQUhaINrMAACnthzQljADuSc4JL/2mvVNN5xK3QK
6gL/6CA7sDiYv5YDx5mwbESzfnVGZnlO/B/HUh0Oln+R4pZUrmfjww6+N/aJ0LH/yssNz+S13fmp
etKuXAsaLe0YMdXuuGWR1xId+uIof2cHF7BKL3IY21rXHiUYyRFOsY3NSpqiR1bQKB8+3ZyFywBX
18KU3w7ASrqp0ZLcJrjtIoAQ8CDl+sxlWldearW43oRxbXamrUJC+NqJJEnlTTS+vE5W1dFWiQbR
xHQG7CqqNXbQJcRbdlOyctMUguF0M/CIXm7KMGCDDpM9/H6HJ2ucGQ6VurwGf7hc237IWKF+MuNZ
v0+QuKdzjHYMO0mc78NlD7jKzKJ1SWM+exaZtfSugCENys0xYhbLbnVDmMV8r3eaB6x+oaB5B7sT
BijPdlS2RBw3dpw7U/09KF4QnC2YMlKZPFuwBV+w7pvm7ZFD3CL7luICrdpL+HWbnsAhfuWgIFZt
k84m6XXCWXbnOB1+r6PHs4PEvZAY5EB7Q9rJgaeqxMnoRvOpa/WWfLigCcfuZY83cQEz8T/Klbq/
zfM4cR47Mc58Tjl0STUgdM/FqDYc0FnpwW86G2HA7myC2iUYUuBVISEjxvKChKDxJR7N90HHNRsp
iMes16AQdf+zFCd0kmP+ZwkFTDUGtVcw+mnqucsRIj8b8VCvtM6IbLC4yiPoYsxRawuZTUZn9ZKA
bXpY1tkq+EKyidJRdjtXR4ejG+tDRSTyc0t0+AehUHAByv1uO5YbpPglJAtuRWn7fgJgIpiqUnCM
0B6LryrM9F1CzyWITSsMPo81U1Gr5VOwIe5Ehsfaq6pG2qrqXMl3xPd3eCNrzpmozCK3D6he2Koa
YNn2pRphcUM60ZU3MHIvRK3X0/vPG/cxhCbOWBGoqRqmemG8jefRLFPWkJXYAKlQ24jVWthS2cQ9
Vdi53crwJk60Dh6aOGy2HVO4PchZFLDCoEQy/eP/yjUgPCbyjQQaQ7rlyWehSIPEjBIXmAQWH65x
2G0T4yOH47BZIqL9aHpBSxgjLjGOtfjKBjglUSFzISgN7iWLD5R8CDdnUbD+qqGQbn/PtwTVywKw
+YNCYZ5DQFreCwB260ek2wiPaw+hMDIt953TyNyicG3fRZrLukYAqJbdo25hDrz3Pbkt33RFZO0B
Rxt315vyQ3FiNhEPmXdYOvzP0drqxUW7PkSSM/C5wJ+qhBHyNrPlJj8hjYpCrFfqkbIiPc89N4e4
htUB6msfqoVxYPInUm/i6s36fQ+QmWn/6RSDdq2BqnWclRjr3nC81aHL06X2Y6DmUeE1BPK1PFwQ
YyK622zW3JaRYd3dYRIW7JOokoDCaWhsFX3aNY6YPYuEifIWQ6cc1N+t0hMGAVRa5UXRiE3euU4D
yPPeG8rNX20EQTlCV0uNLaIXcNXWbHRLA+9ataH5605L017dGZ6lLsyK203EFcJQbu9R8qG3IKP7
NRYaMc/A4B8Fvjg/N/niwAaL88ipzz8xPIqqyTaePUnpc7ni+1w1/zyUH6uew8Vew5/Nvs71nwZa
vSq0iWlflmjon41Iq22VhkMCexPns7jZk4J/VWpe3YeZlyRdOKL1vqNYS4vuYN+6um4VZlkdw55e
MSDXzjHv/5kltIuZXIY4/4III0htbGtYsglElLkEqU12lLswwIKt1jsCYdE0sRZzUckL6cJDIA3L
e7QNoscqun4QJi6oNdxRCfc/CTCizZev519eW1LMwQ+2a0z1Jb4JnIM5kpYSxDkKZ7diM5A5zlhW
iKr9qGPa1+Po0g2V1ZhMjKkS3SeZTSlDCn/GbuwwQBwXsBRWLDrXrEVGDEULor2gBX8zk40tY+kd
+gE06tTifabZ9VDOUlUuSGqlKQaqK1+v0KDFoGdKGmUumn8TRaM8LizGk+ocAvJyODmmIbb2Ch4/
7IXCgRy5kdPdFkLARGzwOZVjKHxm+sK1QIiCS7Q7RhNhMt7YOCPaP0bD2+M6emhflSX+uDWKUC1J
CmZX3j6mrXDX5uJNB6mfiA6YbN6+5DJZBCFLFpFhvCtSBvyVmspt7BM6Ja8x0a7ExvABpfZ2qnt9
cx5WAnj5CFOk2+mOr8UPNGtDTljFiFP0ag85+bt0iRDKtLJ5cGzsrw0X945R3TlE9CMr+qwkLvy9
Jft+taLGDbNzaf5++CuY6s9HD+XpLZ+5lJ71kDlzmjLiRIdPu+3RnLgD4yakxKeEzU4Xx7GVmNtl
e6TgOK4zkznCGsqjOCFLvMTa8VT6Ptz3opGsYfe7IQbBL24BWrnBBxfns3MRYSjqoqlYi7U4p72I
N7nf3e3i2Yes3xUwpT/lgW5YYzgU9FEB4y1Hr+4RJTxqUJrxyS9a6Vc0AsA39fhTeMiRgyP3q9u3
XPlXMeFfWjX9WOS7632niF9w/52G6W6+jr3BsLGMrUMR+a5R/ZDLyJ2K9zjaLDyB4NBOFhK4yMJx
FMYtdnGwvEaKQd99Mlb1cSB2jNW7Ck5R87SYdnrD9SQDpCH94Cm0PzWQfrcgSkNtYzjwbaSjg3vZ
VOmQ2LnotZ7cdKeSnjHbDzMejPE2PdlQyH59JWZ0ElxDtzSqprMOUannkk0SQFulO5lhHdYWI5sA
A+NH77j0MftmPXAdq/Es+KPQ06YYlF52Hy4hVI/RpA53PTQIMv3NdU5eYtZGfr8lX+hpVVwWv+oS
LM0ydqf5um986XuxOACb9GYh2H5mfN+zLs4iGQgLEWZI4KNN4pvTolEG97Y4GrmoFOXMY5QOX5Tk
2OJU63YeFRlkn1FVhcsQapxWGvj2ZLX7jsJ431Ayy9+/9InM2y2P2yTsAOx9+D755pdF9OKOBoKJ
5PDOnHIq8L1uXE9379JxwM678yrIlAZ90Z5LdV8ls+5bBl4bNbSOMclrfAQ7xq3RLgz1XX1Gt8aF
RHpu+P+DzsqLn2cdczj+H75Qw6ZAK4q9lpG+0M+YLiL23gfKGRj6cM1SMCIuKHS+79O6RQvNCSMn
L00HvrxlPKwSwRh4uk03UK4MW2zvANy4RPENAezYBf+WNXdS/Yd0XalXLIvQQN62IKpiyelynYMl
PjoSdiOdYt5ONp2RAnzrELy+1QONQ6GQQoKLQEYtjzTeUc67apuOQexrU9u6Ptt1WwWhsAVgeyiA
+JXmuOTIN+/dteS0oBj0jCNX2+MFcK2+A/Ixh3koZl97oHdIqxLb3+lmzeLfKhmvLKjJqPb9+Qgf
KNBN1oiMfDUl3ltaJjL//DpE+AoVdrcxDLzBjhzKohy9LhM1IpqHX3WKIX4bSrqDuYoV8tNK0Hjw
9fXfQlLqgSjpKV3zWQiKEWNtXyKavB5/lMpRhMTWFXarrFW6cftelA/i8XtxYEGgmVLFB8ysiig9
ig9sR1o91v/RQrMfyM9ICoHGa19d8NQFqJ5vgAOqpYAdMivkZnNGJGt51oRHVz4Y3LJeRXIYrxYI
3WJeYgqFx+1c9F7QKiBZYzKoQsIc1iAsdfsJj01NvL/IcbZBzUj5Ur+mXj+8a18KnqPHQLyYRr4B
MXAavkiv8sy50DxwW8hX4Z/pN93CwNQMUONfmdfOGG0Jo7EUEjLS0XRi1DGQDpPapbvMBsYMfg60
f9fmnZy80l1YNGv3/WbjFjN9xKesNkhgMBGqXHNkUo8ErIz1eN00qO1uEbImPyY7yoOKu4yYMJFG
S5o765tTcBBn7LtpUQHuKbxqT+JvlU5KG56X0WWNfRBefUff2+IVdFMmaOukFxkNvSxSPsfNkWAP
ODf1c4yezaVB5eQPdUZaLYOWVPGZ9EJ7mnYneX0VfMnqs1k5hBowz/pVXpGP3WneKCOrmAonhpwN
q313Ay57FXI244S3RLp/5OXFrUiIsCIko7zDq9MqLrxbdRAW9Z+xmRCmHBd8Q51DUV7c5DSAPTnx
XyxaP98W4lLTMvmaWinJUSrltl+Brzio6SNe6abcSDoBnS+TVvunjSohT+jXB0T2NamNl05kPMD4
tU1UJyg4wV+HTh0Y/8cD6o+EPZHNFEZ5qxcsrlkbDb4FweII1qntCcG2GO7RtcC9so3iP4ejowmd
itKbo8QYJ2Xrd5qQuW8DGIliqIaWpFfvwUrU5e7vb0PlqeI/0NDelOEIV+60YmhtNgz9u4eplJ8l
MSS54l7sHYiuYUal8OC9SySUz5GOJ+qTPdVEfQU3LiZYeKtrn29qR0/O2jMxYBlB8em/O3R83kVs
4q0b+0cCCuh8WN06KgQERo69mbfhHGIPt+al92Ws6s86dmBTrVBpcGRcbtVXOsJ++7EKRAK/bWbn
EQm934jbUpFkVUxuGt4rTCzTmgij38dINayLOab+N1GdXYChx785wn60uk6d05TTCM+KDdHaKRs3
VDDYY30Y+wkC6GVUdHmRxOa73ss88sampxvVdbL8kjY797u/h8WLJ/mSmjK21EVNDH/9Sv/nSTTv
Ae6j+dmYlffHSf2l4HQj789IbIFQdoykKccdzfQutt/Pz9BkYXjr6UGMz8zz7iyZymnf7lfXgst+
M4aJZbTjfpHPnwkLn4a/MeCBNHwsF+N8NBBepFNl0GwWPqhAQMgUa8v8VNrQxUq7WLx2iKS6g3BA
MXH3xpLkWkO+ewMtOwBrr6yDWfB2hmG/FzJ1FvQho9gtECp4cRy3sByK5h4N5LrCJsG5t1bvQamV
m7WR1m36imc+8FIEcZBBaSJRjulHcZEtzPpNOjXpLyKCwyWvyBUnGSASJOfXuuQE3i9ZjCbt+nXD
3CXdzhHHCC2ZbI0YixKuoVo3WicY+4EEL2bKhPdq8pp1/hPS8hjWwIYWBwChK6YR9l9KY/SvnJnI
TmNEDwsT3gxkI/kcHDWYuKMSbmKU62pAUXTIl/zvCwbtS4FfEDbeWdFpa/OtfztXXvj9jZCNKdY9
F5/AWmbr47476oQ4AnwGyDVGa+KyVMQ7YPEUd2m8vnP1p4V3/qOoQ7KQ2cdocTXb59exjKbkjJgl
+l2Tp5vg89jFxbxWVfGTiJBu0yrvSpJG01B6Q9y1rWYe8u8Qb6hmNQrprrzlttWKgs5Fb2wIK8Sd
uWUaZ3KSVc8RyiOWcsvMUzE/BYGz8On74RHJr39V2wZZPBL6kNyAKa43sM04Wx93F1bvkNkTseJ9
4nhehjOafCVdQGP+s9Ja4lWbR6UaHuXUyeVROPGRic+nGXvitf553ZGEM0kfkZfz319tBB7Qxd7q
mljTika3+guj+dxL6m1v7ELtTCeuE7qSY7Hw38IJmVVHgp0rQQUgem6joW9dgyvBwkkPvx9FieM5
T7fTNy+TbmD4vRoWa++yiDxb0N4L/Zopqe2WVJBESx/cIpO8L+91dupt8XKQbSd4sQRWW5dsoG9t
RW7a1wObdJdoB1q94XHmZZQIS/FGtHBm93vD3/Iz3w4iDsp7JkLC5xAbBFUgsNF5oYL0wL1nJfsn
1e8BnhNuFTPwk12cEcCgUnrhKTHIwgLyF50a+4/xFhYWLvq5GaZ6o8e3HWLSw/78qum/2Vem8/VR
8BGHZsEGwmv/2t/INkvzO2/kZph/ek2Z23ch+i0UkvKu8LJ+I8y7YnMA9QEKQHKv0wYMGkQxWmVV
qiK0QCr6qXynyH5MyGgc2V07dPn7RO1988afZToYt08CqzTMMcWJ6hEe/DTtcEg1NSDaLgsRd3kP
Mn2i5y3+8wsxPNTsbvFWhP/PsGX0zB3xQYNOdX2pEzWQ/zWvextQjinUU5gBVmiXvdHxCO+zCF8k
86EouQBfaaz/bpidSTUh6pF87RvO1MJ/RTtQ41DhJwlEvnYTXgMwwObMMfaSx9NZdYQnX4dQLxqB
srNMx9XLmiVV5ssnOd+eLjazvKInkOApTtLvo8Q2r8KF0/Gacop9LpV/4s+uya4/DOF0jMBuC1b5
s7Wqw3WlSHO9Gd+tCdBYE4g85pOZCMKmKTirjJCd4dLP+rEx8csg54SIHcARLoHZJpJpK6UuXu/i
aeboDSRcBDnuMdTxCg4clRtPG0nFvCf0QgVTE5Appw1T/Lv1Y61bXp3oM1g7Oc9qKEL+49PFfGV4
pwsmmHovT7M0lWnSpFjpTuqU21aWnJA/61R/Bv3L1j40JJZTUMMYaJ2PrLygjstx7kgR+XvMClbW
avRX80JrKUlQUYu0/Pbc3I6WZXj/BJRt4YNLPHZAO/QkiCjDdYBjYfd3Ce9x8uZ0kCHkTgtJiGJH
OM+bp2+NS3rdZ0G/gnt1T4+rcJXKojiUBbbi7AOhJsZ/UqJoi1KC81ZAlbX52Pt3+6NHmv924onc
EIcH/bEYyQMVFcKoJfAAcacSFDqckYqTRkPOd8bKe6YEXa+LeF5VASfcVT8JdY+qEscJEoNs5B93
Mj20yP4cYgyoQicClxMlPgrdNefgqd5kmR8NDewntNTS4Y8FOKazYM8za+sGJOKgHs64lFzMPtZW
E815cgJjmVOAX160o2UGumEgAvTydLcad7JBX+90813cT781jz4ZFsElcr+Q5F+3vReGbX1dc08Y
eUH0fD+skVx9rYPrqff1hri0yoExMcG/1esP60W20ldGL4ARTNHtQaJVrFhJvJKOqcR+jNYJeKbS
Hz553Mpptp4s9+y5nTOeSZlwMQss3W0x8+2UYKFIb4hHbirLE4dMOQuW7X6Wr0YiV1TnB1zdNdEp
U9EILg2dV2UMLxspiXgujrEQw1b5QD1Civ2VlQ2Nc8MviZHj8Mg/Sjd0rwrvXpWL4EV2hzCZ6tUg
kKpM2IWdD2EQTal6LRxV/EGZrdczgUOA4G1kwQJo8ONuyiXxawYeZrOQGjY2rSHxwynXxgJypp7m
MDr93FwQwooFoacLCQKNfIFP29DsRcATxwEod0Ws6NBCGlrEeG4+JTAF62tg10BM+60jbRsgY2W7
1s4kumLh1dbX1twLwnw9XhyVLm08KX21AZ8xW8uq8ZnvRow9R0KJPhcTHcUllGVmO4cD1rg7LYXn
FpTrA+gBB4jnPNrw+slen/jEkdOtLjb6+8sATKh3j8ieECkJ2X2guNkgkH5mCJQ8t9xZUte+A+0I
9A/5wjhqHl/huXAwLwOt00Nws84r/E09WN8C4hdhBr9eT5GsWJHoDXKdsvIsnTFPuEEZdDdS3H1V
rU2YPvoEXxXNxCzxudmMtVPqo54fkrVr9F6w6P10FiVLmjOAmg/bVleB7Invmkls8io5D/dTdvxK
I0ylOiME8O957C2n6fi/RaqehycjX1K/HRUo9+x2chfX9KBJnpl0zTmhf7ZBFmy90pAJ/VMhaLQ4
zGLjtpUHkNIYuH31bgoMtyXoeL6kGpcVXBLzExko19KmTl6V7+xg2TTBBa5v0+AqMDFn+0s9iFa7
SlflD/+3zGqQhB0Dz1lbhyrp6bFfMpjqBmcvoZe98F7k8XkycnoE63llKKGwNj2x4XJdPBHP9eFO
fah3Ig42g2kBE81H2RiIYPWlwy1C15BfNORkgfoEl4scltzCRdm+LVoBgAoMj4RNufXqCyQpfY94
C1WLnAiH6vyv8+6P5jWKba3Xiprmz1/Jdb9o7WwViUDBtnnHEx9eWz+9opfOhlnZ7t13TCM/AaUl
3HfhQA0DSG9QJvhTFgXQJ2sNRljyL0KcJs67ql5FFoN2JGStl338y01Anz2ZAz0QQHonxnmfS02n
ft5tmG/I+hMIv8RUq58Gn9ngZTa3nGshFcfi1e/4g0HAq41m3IZt9HTGhHKsunLjwDHpvk+ACGvh
H6iiyWQmmqD+Lk8l3/wNJEe686jzrNU5f9PdWxjdPG9kDbSNle9VJaqCrCopdqukVbl2+Wko3UgK
0U3R179KYUe0cNro0zlyXX+R5nk+BJI8BRasMAOO3LaZy8C82WcJd+EJF+Zn0A+8Y1ke7R8lqRQy
UZw4TGNSRMgpeYT0+GLZnfrr3Sgokcv/oVHahRMoIL/FnP8HC+0HBmw5BgGfD5GzsFx0ZPEPknib
bM3KjuKwAGMjObDyR0pmq3nWBgYDkPokyryXKOvpJ01rBeFmE+uP/YwM5GsecXVy+pgoSXStsg/g
ezgEFBgTnvROEof+Kz+XNpoHNCw5xMJVP6QO7TspVpgUqvbdwuAarCoVqBPk5cnEO5ySya9wW7j+
eYRTdC+TSM4fec4klaWlTg6E88pzrgKu/TVr4rrt8HaPbcAFyNt+kHSFyIpKxTJ8bd4gzNchtZ8t
a3n+VJPMGmZyboMzZyi8gbrUv2CJ2DVAuDzLnA9y5/ryGkC3lnvbl+JWlRhJw0i1M0NIsMOfMUa+
b3DuUmn+uh3HCJu4xgvW5bqlmFJkhB4ZiaJ0diW80XCd1Hr3giQcyiW416K/4/xqA/Abw/L1ViJO
7lEweuItcA9O/mFVxdhlDvHB9Q6Mr4scKAaiqy/geR79L0OwUOSCHUcL7W0+9kZViVmQoczdm/C9
kInkxjIjZl3G+2DTH2L0cnUaTMEwErc4dmqbPxkS4xY0nwG/X8khwb7N51vEbq7Puq5qLgzbQlf/
15giWydjztwR7iA/eAJiMob3FYjCtPaCp5KjiqZQKnguE+zOgG1quN7dSxXolr6wT+rJFs/dexpI
9BOo6Gr/wBiQ8xgQd8/ryyffB9CaXoar8vR+K0VDN04LLO39XNJgZR5djz7MTzHl7tfBMyvjU4dU
ijMN2m12mvIcnpO0TMpqvsmnx70wpEkXR2CJomMHIhVq1V5uGu+WPkmw1yTQQhMBOPMR8QfROvku
oNeVPyZ/OhpoYrNrALjddYyMmwBR/AlygX1OTJujlhF/SGcQ72CgU6f6UYOFVo0+fCGjV+Cjt7X1
pW/3q+tZBeghGomRVJJpaSpjf8bfovjkHQD5nE2ObnnMP81I/kqu/B2EZHkIdZ09fyb0p9Dc2VqK
mKynk7mBfZ0B3ikgzKaEampKbLr7Wu+bFC2yBdCoPjBlEwHU+AWyDsOYKmTVUJXAqfvEWMsj5dN+
ySshd8sVGFjqtNz12yDvrMOtobzAXKYne24torC+uthxMHR5fkSpH4Rn8j0xJ7CON28A3PFg+LSS
QzVbcS5xYk8Mg7nKqZME/hVSPyJh3uh7P15TCm7xQv/0Q9A5Uy/W/ZtV7Z2L2DBa233eb8cON0BE
QDTRmoMTD2s/NeFg16NWvwM3MESOhwMcKEbOfc4FIsdT23rAUzEVF2AA99+Wpi9+sB9fGVmbwFoc
pbEu3VIvPv1I0WneCNxAWDnKqRSjElizG9cOWnoRdh8gyJ0Rtzz3hal8+pFT/v6vSdwwfpGnHY6W
gxUApykRLwboSdiGD4vaj5vrq9hprmP0qSWgkI4hCSX9CQmhJl+/zDfQJ3IuIALwjuh9n+0uzIBW
qEmEwrrZ/sID5fZ1lRD/GmZ2wKCSbpArAqYXA7e4N8zLE3YQhfVQT/ECoTCAv0UWLxURlpOub5iG
4U/H28TfDdKm+wld9PHaHMQrNfy+9dxRBjF01uGLrxPOywbpjAc02H8t6lcoxeNFaDYndH9sUVsX
PonsDMNLuFLsx34t3S+l2lsrGH86ZHdHvDgIkqHkAtZyYcQa0oy6m3CfnCRu1Pe8jg9kJo5MIoXE
BilYMzDuL0BsUyLE9wkaF8BUw1Te39tfzQ9ddW/gytp0RmWsrzTCWsrGHMAEIH8C25kjPMtAgZgp
OCdV7hmdAiqr9mxS2VOILVvYb+Qd3X9g2ZOorf86Jcl4K9o24s7ZLua8uMYW5pGWIOOmp/V5ygUg
U11q3t/jvZ9ZjrSlN0J12CogViWPkwQ2fB/6m0CPq+NrFD88Bh1vTZRSJbu8fuDz31pt48HYked2
f1B6GRXLvJSQxibfvy8Pap9kSLhKHLE8Mfv9HkuEN8TaTVfy0q3MjH/hlfLCG3+nlHa5hNnuZQhL
DYIATJlDVfvaipKPatMUxJ+htgiLb/lC05FHztJJJ/7w8N4tM5l4IXo7eZ4BA4UKF2FeIAAy4PBB
6iBlhYHB8e+hbQe9lwJdlTDfpgU5CZl2ADCKxUakwW63qLqCCx/3YCYkHH1RT1pno42GLCwJVoQ6
etDrNrSAUSCRZM6GePrbxuuCMktHXkRexaEr6TJxUxxTHGpT4xKvHqd+o3wWUBb6QLU1oyRIIdzt
gv8dW2skkrwQujNJlpGNalRr6biRrJtFoWTXY5Ll4Gt4Fy2zNcVo9OUyM2d5GSGXqhXvNJXk5G7M
+z4xvocsybwXCNcbC92WqSsfro3yHIg82LlHmqaBuzUKE6Np4t0epW16qHLuJmoPpliQCWwSJ9Dd
uxJby1SBEI+avzOQ7gf7tVa3eXUfUGW+oEL5o5HBnbbC5Rl1Ha7AAInhxVtp2A6ghWBd3LtBbZhm
1KBjsFaDzxPg0vZuXwtTAP1bY39KZa2aWKlDs11E1v9ieK/I7acqZPgEtkEIhCvscSBw/eQ0FK1d
25Uv2WirDu/tl3kkOvc15PTIQqDvuh+eNkXmny+xeXW4R1zrnRcg4M7You8yGmtYajp3zSXPrUGl
YJmSTa3xJNzP14MSnG/vJ6C4bMs3+9ck9m7fGfT1IAHt2WLQeQsPv/nBzfcaapfHYUlyHMf807KT
WhokVLBlCgA47depOyXDLtdg5Wq2hTHrx+bkUK4ieVeOg4eAXfFOOYCXhi3lNJ3o1f2Y21lb0jxP
QAxWVoJKFAYOLCEixDQ3cRYLe2+l9OOVOTEq2OS4Nd7yFtWVZXHQzJbB1C5NhvQFNiY/LUGCEUDV
PDTxbi2A7Y2g6qIJsN3UYtFF7GUJLf60C2s8/ZRAhqFuUWsHhjNIGC36HCFse14mX2TcWN2h2p2L
8GbsoI/2f8J1LAgVtOckKjb9tvnq6fEtEVcpNXkgKP2yuQ/1J17Gdm1Bd5Ybx4AHo8mx+Gbbw50/
yZCNN3zLDgrj65bdPcgUgP3uAC7oLiVuuUA8z9RQ1lsLse15ZTtFoFbujgnbIzKZPPbDmmMC9g3c
uRnsiAIrWcvFg3zgGCOD6YHmG+gcuobNXobHEElw6fGjI4iv+UC8TtmvXNrJQmpIOb3WjlnSzvJ9
5c3879CrD3eYl3A9E4tOKI1S71w8GNRdYF7xs8cp7AD+nTzWV87FoI+BmmWqUrx/f7nx7e7NG+Ab
2CtSLTpPAvD3oYHEJ7Qf0j26BDeJlX27BwDVLPd8kMyPd/J4xVZIrkuhW1R/UO18kCfK+OUgCDjJ
S5kMklUC11RW9QPzERs9to1lGi2mmi7ONWaZ2nqiMLK9hiLETq+N+CEyHVlNK5wiQpEc+Soul12h
UsEwPQ6iCtpVsJnZJTPlRb3FwN4/cSbFlohstHwll9q4XblHoCPKVVlqNlxCvf0dp8ToLrZ57zSv
B0v58bUw9C53ELsglbc9/bbB+KJLzn/HLrBugpa8mFMNZzw4mGj1PtQZ+3Q86RzH8PJICdItgzgx
5GnBHkqyj3/pbeP0qJs6VmaY27X1E4qxT9ch9XyaeftS5sJb9tBzHHMITy3XLImDx2kCb3pM/Riz
Kk1ydX7NOIhEf1DegvfUWsV9lK75tOuUmm74ruZ2fM52MwOhGtsePeepQMHLctKoS76H0PzqOG95
NPVVZBMLIktPb+P9PVx06ArPSYKAozzOZ0k9y/FdtO7Sy0T1Gp/XHm8zqdH391skVyd0mg61R8Bz
3m0apRCdPnPgPQIxvc91/DA77O9MR+g7V4iLmBF7qqpd6uX1Jd4j4Mza4/owY7H9EWjz5uzSB5kE
cGWXopsyMiIq4pB+JPYcOKxJfMulblhdjeaYMGXz6XPDyDLLnIOECIWAvsHaN9AQbjPqG9k2VcbR
QaYSKItDVK5QETRsub6x4e/4rCa1S605KbfADbYjmIA+4ACp5UaKUvpbJDE70LtQDDw9juVHm2BP
xIjOafjo181hXWZ15zQXdPsCFr9UTPXKvvHcrczVGFREiTWoCOC+XKt0wKOuGeNK2w1v5fVH/WNh
l0vGTFs3gE8DYDS31onXyTyGUDbNnDAhRMnXgalGs0k5FD4qUnRHw6CtfUQrQ6Jn0DIf9TRqHOWg
+SmzcMsPNoQLyFX3n6w5Efk5EdJ09dvfFOgMe7QeXlERUSr9DAuAsh5p9Ht7Lw1uvaB6PN4GBP+d
Fvtil+HQcq6Y/TEalEuZR+4CwmsK2QE9k0H/QmjFjzu0o2yJlJv8Vlv/9daJZA75+W+LTrODlM8H
7pRiL1UT+vEOaR31M/Av30TC6i/6SdtluwXuvCC8SDyvpbejhPxUQoDePt08k1hXXA6PgVEtY5MQ
IHd9iG2r8xXCEVlG4xWPzDfMsTz0C7Nh0FQu9dLgQ5oyUPT1PfP7jH/+UDxaIl4XfbqzqooSaU1+
dM9dpKh0cVY0p3yeoSvPlqUdT6qXXTUqA8rqdzvchlPZruJtW/i2I8H4yyZuMBhlH9++FVP/xgbb
z9URTmpFqrcyvEsAWFXIRRHSkNRbqFlbbeaAvSSKEDGc/l8mkQC9LmLcnNTjixrNHCS8PbmChLyZ
IFOagRB5kNaUKHWXLXfjAe1rsqXLerKM0vNDiRA/pFAfwrproAVbn4MrSSYJ8Sr3K2cqNcm+wLXs
4xCLDWa7bqisTZjQzYKbFbC4+4RZlpSQJH9m0BCv5EnWFAqTq3hFyK7xo6Ty2Hp/iEJ34kLH/kAl
NE7+UTOapwCU3TOzlkm0ZN1rItG3c8guLMiss+dn6yNWsmCeP8cwz4o1XUb70cltCN3yKRcvYcMo
oGpRKC7tqPFwGcxgg4tL5h3DaujB1QdlNibGOS/WrmSfgQ05z64h5TOrklOEb06K1IhnhvlNHbHn
PHFJsJRbBBvTQ71izz3tl14ZwaDKPL4XBDxLbhz5GzZlvbzZCy8qFb74Lbx3sCq8XsGymO1ef8wq
QN96LU5RFwsY3yqa0/htcEoCkPaW6QmW9BRPNM5YnzZTp9rJiPbPqcTpk9nwWW3Li+c8DOg4t5q9
iaoE8oxZWVJ1X9Vd9zZOHGnuuToQS/ONmi00HLwUCsb9153Ew/NXgXNPYZNL3bQa0+W5pUoyUgtp
Bf2kUi2asjiQodRQAgzg0zCSS2jzyhKzQNo2NWz1LGWZVBz5lC5Rz3bsKYxr/i3W/FqWGxC4sgpg
5Og2qoiqqzW4SFfqykaaIoPQNxhKQ/UveGFRsT+vZFyu45c8kx46D5i4A7LtvAjwF7ICT9zOThfr
DpvRa2qBsc6drlPqOs52JQXopKQNk6hEIp6UeNHqkmt5ucqFRfhAyTVAvY3Mf0TWYcUTcnAKAOSG
W17EOprUuBiJnsTHY6p7FtetT9CUHz8ffjQj6s0Cn5LCkavwyIs/5KMtR5Z8W9oWYv1EwthFL4BI
RISfdQrDrxtkLjH42sq8Q+K44PpQiHokG100N2cvboqDW0+bpHiqsu/jTEj9XIdG+nF3/BqvVzdd
QP6998FUh2usV2KDc2gdhAR50H0yM9wMJUWc6rMfxusZimnl7fM3ds7guJZdIdpwbESl25dW1wRA
byHNhZ37vx2x16pMflWypTr/URj6F1s82Q/RDxtYEFYo3e6Cacyo6lwILx9G+/IZzXHsRr5z5TSY
JUEztZFWdAoTb8P8nCCRj476weQrRrRVMW/tqB1fQyBwx86ZR/eSKiAVwqXqH/e7faK3nb3hRDWz
zRgGs7c0Eze6hiXtJc6AfRegRk+M06nxruwAQdNOYbEoXsf/4NIoiORu9+YMBGzEGY1hwyjvpl/u
Rd5hb/6mmJEiklcrNqfJ/zb5EIGoFkjjjdn8grwS0/ccxxGES9eRBnVkPTKgaO12mpUV0CM51hrR
dZK729jkGtR3gWwkD1v4F22U8uEgl0107w2m/VllZ2EZkDZR8Pr+C1Kah+UEcbHzHPfvJRlXKjWh
GqpPmrv0FvDby92InZkRxe8vFDQzPDyF/5e+kqVUp1xe4o8vuscHK9vRxRtULN2ljEXAVL4jJmqC
pH2kh0JhLEGe+vzr0rm1ujUxDiD7N3JfgbU9Iz3b9LaWrBQEUrGGTsP7RzSmPM7RDsaUIvlR8I+r
SeJC5flsAJWuuhg7YxMbst+nIuWgOfc83/B8+Q65b51oLB31Ynu5DIpGipmUfrl224mt6AYoym7/
m14gwmkBCHFrTmh09mFkWYHq8ikkTJeEe6P+ZdbHegOdkMz5nhd+C8B485u0CnXEZ7pGb33ihP4U
nC3hxJtWMStB6UTXGor6tRrV6QQYXeKo+vDdT8ywh7A1BIpytBCpXKekL+qohi1pVfAFO52ayB3o
Q+VSRgHQGvDOpiY+10V/NvhBhpszT4kKlIZeLUnMY7F5WN2ItJDaZ/FVb2YQL+AVx8586oHwD1C8
A2ckkrkqye1FDBeRx/82TzTVroJA2Qbfc9fEgV8wU5alG2+AXHqzLC9XaJI05f/sMQeldC7XDQLf
zumI4ARQT7J+WbLQmGqBBxmBej0Tkp1uGsVKZU129thbplU9oZL1Udp4glQ+9uqm/wKoKZHMiBNA
FrZm02CXIA1Gso0kOmOgLgAzJ/nJSjcvgyjUW7AOtB6+Ztd/di5Apcp9D1AFfVc6Tx31eaFUCG2v
gIkS5VK9mBHq1rPnZ8xpAKBQY+hGhHxvID8TzPmh7IorO5Xn8tzJMeP1HxyyhjybXYPvVKhz1Guj
IHNmaB7xxypjG1m66sESdYvXiC8VfT/CLoDXJcVSyBNxzncnivlKucHe4FPxCzGXg+HUllslelpJ
XlTABYC8xaPQP4Vn6RKm2HmRe0ipzERkGJi5h1x6cvJQeR8AFkiniCyYuarGCJig0JIrDzAIpWuq
ZyJ1nh9Mhb85P5bFKvYYAodIToWrnvr+fBZb+jIZKjfNEuh0/jdJgQKdBScTVFihvL2Grs1yqTv6
nCRqISQf3hwsxA+4Fd6zzxHeJCL9ponxCY0ZLERXCsp8F64pk9/XhY0TBsXEdbqo/3nNVe++wqyA
ihcPLSSTO6kEZEcH+aVv4Wl/n84aGCO6x501MmYytfY4wZBN5L90alfzMOWcW684mAShqTwC7FKJ
KSyPny/AZ9+/co5Guv+T1xH3DzRrtPu8AMOiBOmLL3OV3dGkMPBNeLtjvamsxQxtInCOp6hhX/gZ
bH35wIKeGqycKkCcaZdMVVANCpOrXWAujfufeJf2PSULVeLE8lLleDcy5gFq65NdhmB/f3Y42WWn
+jMHjxcrl8MpO9i/PDLGomA0C/QStlg1rtMPiy3DD0lZbW2bB0d0/bM+NqVFeP4d4Sv51jdAVEA7
B1OVR94OQaHAaWpQVrUT3d7qsqhupTqiWQ/n7FBqr8GGJT2vFg5+SlkP+XJYJIa5i3YBXtZ4QiWP
bL2bxSRyeZUYk087Rcq76ZzWVcOud0MiXkJqSW80+wpalXQjFE1rMX4XZgFZE/WhWocX3xBOKikP
t8JVMzm1UKSPWZtq1J1YFWRLzHEjcrdiMd4H76YoXkhG3kliWYIUmjQ07+/EJ9A9EzoqARj4BFNe
ML26Wfs+UDoyLApE+n5KJT9jTehk4CnLtBImjewzENZdXzxYjpM6SP9R2AZ+XaOPHXzMoh6dA0mg
B5Q476W8W4syXb3s/HV99ZSfT8FQnHLDi7shjgwfbsLkrhexa4kPDloCbiu4ZaKymzh3viuHrVi9
Htvzla4cpaxKvtKxvP0tAORCpVVRP4wsb1Wnp7vc4iChELcGFF4P/AlA/00iwVsTr4ShaNTamQeW
bqwcmP51EnDvtmgrFEnAdwUfLKsQP+Mh6lRWJYQGle0dkdLyLC9UO8J74NShFTISjIUJ4jdH5s+c
TtFJlbZc8UbsVS2VQi++Lroj6p3i7cp3Z2oMN30mXGOLVEdJguAvOYRlrhqxUnbOmYv9WA7HBC4l
7r2jEQaZpzP4JJl8mDEdyLLeYwtlcYS9K8MDSW0xkbovuO5mHXa6ZDeMnqCmcsvcarJBKd1XQJfa
g73T1fOTHXeQXsbuFc2/mtYasRPzq1Iwd+rrLI6pmFHeHJs/JR/kOX124RM+VuFoVPZSsUS4APgZ
yDcfMWpajAUoCQIPaXucrk2DRBUGDsZ16MQ27QFV+B3CtlaiRRxk6NlaEpSX5+FLFtoi5dMDz6YX
0QLflM0/aPahsjeiJg4433AGV9aUyqbGq/KGaCBlQZsr6/MrZNVh0cZoRuCEu5z3LhwAfiK/9qKC
xnSDXRgkCHKgtEfyVHAtR55GdCboiAzAc51Wtm6U5k8LfFl5TRJRcjBBcdQwlL61B/iDuuQPDEMQ
GTsWS3iNGOv+vSgjwqSp5PZTLRk+y9au4nzgEwsxDgD5qj1/Nbb9XQUEHAJi9SDk4Hl5UBzLVwOZ
opysh9snrKm14yVUcw/7w0OhjAt3Aw3Lkr6cRqzOZg9Ocg1VAY39T4R3Y2X6kEVn1De+RcxW7KiR
xvfNo+SLdy0T/T+qKdQI2yZ6IXsy8en4EZ0K62Qkh2ETEmKhDpaxVfydQ6Sf9nET7KUVe9uW8y19
7ZrOk+k+gd6qr+wHP2VN64d5F7P8wAvZjtQwzX8vRgURfe6wP/O2TUWwouj12jISQZPcn28slG87
oRmzECeX6ruOM9N9mZsQ+SN/hnP2DfPTVJefcOgf6YM90SWu66Wdv6d2wRODQrUdx6EcrdLGCF7/
ZQ/kZpDpV9AuMKt3ySu1AJEOjAfqiLbq82VXW/SC341wW/2BQfunD8VkacuQCLTXJh8ES16LptT7
nqMTOpXGya8T51zE0FjjGtn9SDCCC37/27Q/fpxOCc5tVHQ/h6o7Wi6G3TiQRrRzvyUw3H3t0pre
gsvCwSjpUIrjASHfc4ssPrP4bu0pt13NgUIbckButMLYkGkCILi2FYNl8+bWVfa3Dv0KXBpHLhAu
CNkE+mM6Q0KsFfWZvuGhLQhegDz1ULxfuZzGs1aXG+kl9sPfZPKw+Pu0ktGLtnDbGg2cKGxdIOyH
7LLA2mP9aZyZf735YnVwOBeFHbK3aMAK01d6duRjcSG/k8kpx/S+ZWvzSw6PgfKWfYERPphxzT4b
Ri/UgDwK9/tvRqWdsNLlXwYEh1n7Op/EGoeD3rlX/U0ZrC2YC/G/nIc9zPaOjg6eUKjFVBVNBiwb
sHlp8eN26t98I2HROjAKn0i+cr9Vml2pdnb5cSpeFPhpOwr4eRCTPyCtfkb+wt9bwvxcPAwbNGMA
HTZ2LkVYtJmhA8eMRKnAA0QBl2g1vHqVeDLyLIHPsw0TCJmkA4X+y9ac1jQDn2+JQhlHgMHRak7D
idcCjijZ5elIsyLyPuTx/N4QIdTnHxNpMTn+HL1RikIQle3WTpC1O3cyeuhlAM+4EggCBTywMSxz
aKKndqApkI9vd2F60qyXGjvEyNYcIY8jGk8gr8kxsPz676szgWN2VHfJpfFLTpkAkxLyyKnxL8q2
L320Uh5tw9Nkh8gVSWFrP36Q4PfeHkKvOwIsTPZyORzexdCCnqPK/w3D2Q6jUo0SELyxgQMs2uFl
8Wgr5mAObFFEKa9p1Tz4RvprN85dziH8Pw0Fyhsztycdf6qAOkcREOkHlLKevEB7W4l+il/R+ytR
8Q0hJMH5yJYSfXZRv5MaFItG8cFqrAEsRrrxEMSl6IrvPcJljgN8vVqRmyjjU3Uo59FE0YMp2IGr
BU35+1ZBVLsuQKrXPzPn6pypPAI7EPZ2SE9wGiaqdDWD9svcw+qdypwdTQO036bA+GuUvf15JnM+
KLmnSW6ZXW4FnAAQltjflR4a2gsJ00tBX1+/fgUBKYN1ouPpKdBV0SpEOCA7ROMCMEMTmYnomFps
SkAQqQLYvJFVPx1QX8GryvTt2lXaGbfWJZqMm0S/VUv9vzDIhOiRG+GsLUdzcBtmLUTc07/4jKEy
GlPWQK7R0+7GRkmW9HUP1fJTWdx4K1gCelBRPFNV+9ypTmYZASvNcKJDiH1RIKUjktySixoG77hY
IUpSe09Lk9aGp1iceAjGs3vC8teBa56F0LnIphTFbQhUBk9lwRGSjDAAE8LNANAJUbLb1FVTU3Ii
vRw5xQHLvxAYCFt0sK2C7GsaPiycoHhRpsZv9J46pvLUNNKB8ZyGfBp6NUMsPcA1hKVawP5jeaGH
XtliegBOjYt22md+Lsr5kbWvNF8ETRwUS02Pnq4dxhgvuKKp8szUcI2XIMT2H4eUluI8PJSLBAfN
9JiEWgitA4rhQkCelXTpqifVhaUoPlQ9ip4Q0IrswUg25qovf/Jq6cdBGXR6l5e4qQKOCAFja6tQ
k1cnAHnD7zpcJXcRaWUAzkJ/RgYvq9qikTpAOAiDYxKAvpwKB4G2CzYdUdru8+9a1ye9CZx7Pgy1
t0nTWr2uzXjrVssQ4chN/9mFcWjYfLfvz2GvgF7K8lLNpz4AVu3vd/KOvX1TIBXHeMNxgq66CS4Q
rNUm8CqeFhSShaQTQdRIhb92pE3gpCKf6j1eC21IB1QaL0BGptWJi0D3hasA6q2Zvv0fM6FBoQoF
BmIsCmZIjkPQougHFk7Xx4AylEdEqDffSLhmZrKf0RklEYjoftZj6rvw5xrfHJHJr5RmVevs71o/
xT7dCuATNZEyu0BTi70Kt9EYfMV23bE5pq2YRX1xJBWsH5xQCPfsVRrOTGtQ6B8YeO1wZPT5dcHl
Kd6CGQjAfA+srLjCDcNHHzKQJlSqnVthtCT9sXJJji4H1orDxpJkiLNdl5FawKAn6CHKl0Muytgf
TNkv4rqoaL4PgcILQvNKa4NGlHrhjXFluCd+0iRFvM4oysB0fIiq2q9SAZUKMwT8xbRvq3+G9znr
TrB+Hi3L4/jQ+nO20sXIXhxLTtImh6m1C/hHW+C1tIwTgWr934w+Dk+4Ncl74wBnYwH2zH8mz2fE
3tqUwq7ghEFzYpA1mV0fQYUE4onZO2I9z5XHpCtsiIbYU45lfeaZKIqwjojsv6MAk1rS/ANgsic2
H3hTmhxItBARHfnoSckbnierIp7jONPpYg57/CYttIK4PbV8ztJwydRbugfu0pX0d8J0DdCsCkUA
ZK7gN8C+SEehB8quYTfJBAnyCEV7+NkYPO6j3/NbbxTJsCNnCj5lKp69Op6iOEWq6qwueSu480ET
QknLf0tk8qCi16X2QqO4e1xCS8I/8ZPlVXp32X7AFRrofaWEoYCsM/JkJ/01WBurZ404FYEkL+I0
eQZBkRcdZiobv3gRrD3SgqN+zuwAR65eQlM2nMSisBCjevoXHUspYyW9CEFyyX5iU1h1qTCJykqw
7PWDWi3HufcQbefgZEIhb/0M9kpUqxUmxaL9NaMb1LrgQEEN6Chr7Ccxh5oP0uKM1Lfg99ThtglB
y32AvosagX+8g22E8OQNtDmydhDkO7iwOC5IYHcpzT2yD6gH5scLQ973mXPKTV+ZOkW8/+jM27Lx
tZvYRJer6Vk6/DV7bMHW6amQPe5gHEux6o56XcEK3TLsmnzRLAHSoh6+f/YRch5Ur3rVYvOem9Ql
WN8uaoHc21lTlbKLhj09zoESCp7vVOuD/YomFAlVEmfp4EF4/OfOGVJyqw3K8t0oXVLFOBb6Cf9X
4M5zXiAAjFMd7mHhAUnbvg8M3mU4i+MMg65xlpE8RLpBzFBFUEapjTru+lxHmNq7yOsFRaZpgED7
Ej/Uw6nHEh8yfPW2R07mpbm9fm9AruXWgVLmm4x84P84X1qHrcaT69gIaBTjFsIsSlKGA0WuHZe7
k6yVzs0oWqwYuCEaOr8WPB6oiGAsbinjhliPXgIffH4//5qlMWvE86npuAjfnQYVmi6sFi95XZ01
uHQyU5mCiQRocJBX+cMEyh1xHi4AwLibih2t4noq3ozkkBSAKV3xtMJaH5CCKE0jwMbuTxeB6m4h
Ay/oNmfeYozjpAr7NN6a7AzCJsvPDKh+NKyXkkU1gCWTwAESTExU1EsrBlEM6+vWzYogBX5MWKVe
SSwXWGG6GOu4bW3jJ+EdFeFyA9IU5ZvZqlDjDCOdbQm9WrHbPo+8vO/aC3aOF0q/Rd8dEWtpRO7q
fGqQ2uMwfcT28qgpJ3Giq30cbl1yJ689Vg67apcqmpH9cCJ9NvLoZsBI8sAqKFs9jkJ4FVc6pQgM
vDXt1Iy3wP9XyGYr0UVCWs1MLFlYrrIh9IHpG6Qzl45rocVbNR8t2EW8SkpAcMagZ4eItNpHaTBW
8O2cpJjB1r9GY96L6Mpvu8+17Yesr8MvEdhv9GEk7FbzngzLOSWJWmkmvHEDlSqthHv1c1heiXJS
7dPcNJqsJZ4hpQSSjGWThSLVgQEgVCj/x/SyyRH2mw6L5+fELexvg3tCFoDXBkeEc6xS8cTIPqgw
UD8avVIkTYcDJj3/IsfwoydN9HlYqpq/jwFprgBSpXHh19ggbtLFo5qRTjJyOnhNRTCVzE7W+TiX
HHfAUUAeS9HTLPWgVaML1hIQqSd4tfKaSNp3lPDRWpDA8+pfVMbWwl5H4RwIsaXm4tP9pIHkjK4P
+t+TKXp5y/uhWa8w9KfiF02BPnBqH0o0K9j8UF5GU2wjY9RjiGXKS0cZcxDwjVV0SNaRvpTbjKSV
w+UEHImjyg1j+Wx6yoTLeDm1L5OXpa9m4/w08gTDC0LIa5HwQLCy7MCjI0mgBtUW7sgQBNOF4/we
PlFCqy+wVp7X5sKA0FtlW6wiQkQQzJ0bgxsukg8/atS+WYccTqz5bN9xROuHiV6qTjvXY4+7xLZE
hYTcvwFBx28uwZR8cxg/EQ1VmXJMT/JNzimgTFQJF+MFlLZkwlPgxyaeKzIxeP/y10K5iKf2yYa7
z545SwPCaMYQLaBpEDAK9owfybRHH4Q8ihE/QIpnjzPByDOhVu8XtigE5BXFMUxSKcaL22OZMshN
YhZSAV5h1ajMNf+oFLIBnGf4fHCYc8M/FZsTUqi582W+wXH+oE9igZgxepV7aPXpWg0W4E4BR8Vm
2pvtmplO6zz62VwRjB2OtxcBlD85nG/2SCvTGAxD8pE/mvjgPuMlJytKWYi0Rj5gMJ2wMStmFzF5
9rBOeoz3aOs/jXsD6ByCQVlNjd7iMsveaVENdqn+gaCArPObAvVvX/PUc9lo2Y3DkUbpNq7cEppg
iNaVibpFk4zpWbQPIuOOj15yTFEPQeidFTZC17PeJKsLUK2etDS/QMxZvcKMsxvtepTNwx3c1diy
H01fGvnQ88xKgf9uYs7a28k9de8NsyhsiA7Mh0a5EhBVokJa0H4sQcwOd67XDCZXyYfLb/wkvJAW
zzjpqUTsN16vQqNvMLqTB0Lpd1DD1g1bI+ZPM7o1VJyU/Q2W9m4A9tQIK2MKW4ZM/gmAoWYYk9Hg
F5tPKwwnK0mAAu/fgras5owfl6khfuplKSKm++W3Mz7jUMAPvYSU4hOB043sAQ8486mJKEZ9n4VS
hvPRMZmdDNjHZU2eZL8K0oMVGuBtPHzPnd+HLxUms48HBftQfbaZYOvOOklAqUGXe5q60Pu2s90A
dpK3hZ4y9LIyOUQHXvjff0z40+l3zC3q92meDq9nRINBKMQjIJ9O23mqXDPs/HqpE2ipToNDXPuO
Bb4q4OJ58ZE+T8UjuhZI3f8b5ZsMteO82Zgti7Y6eNgXeMn3v8eNazqE6IJfy7sGLC9bsslEyzE9
1d5Xgp5DZ4OWTry1FE+tw6xKO7mmA++mdmatIIVYqyH71At3fowHe6fRnoF3rQx6FjvAuMC4bsWK
lPHkFtA5J0BHlG0pFnW+lYZIex5pzq55MielX/pv44OPQ6YbFhUr9/M4PuPUMuTzdI1XWqiobRRe
UFDouj93eky9wM+s1vHiU1qxjqJiydj/TQIjPrBdezGgpZxJ0DF2rq0wKgoeoOKmKeNpqeIht1tZ
vWC71Rm0zIcMYhKeHX6CjcDKeNDyHmAAr3TFYTsns7jFishrGjx2Xf9/c5angGWriwDF41ksiBEa
zUBde+deSNS2uUtySxYoZr0Zd/lpKhBLwoaqqMrzOf72jZE8qtq0J4AJc8WRvI0N4zVw0Ha5ZzbT
s4rPgKQLXRAOnmrF5u6O2OwF1OjJvDoQD9DO54GW6ve4FaMTxEnKRFbMvGwfXRsjIsHBjpqz8OJt
MjD/lF7/FaT+F3RIOVzx4YkJWGz0M9/IfU+lO925sc4QuO8UgnZdHqCABg6d/Yx93KkHrIb6qyE/
tT9CnZwLuq7BlJoJypJQkN32D366web+UDKEtoQoN4sdAVYxSE2zrXSioxNdYK4bu4Nsw6JJgSxh
aDfb5Qygf1z1jz75ZKbu3LVNmwGUJ9HIoxTzr6VZEUZBfV5tpc1tMt1zDp5jmh8s/9xszx7UtdHz
W7qdxp9GIzxbS0GW+5kzTPSliTmE7KyqhnNUbm1F9CDNll1wnOqXMDKhiMc/VcZ3/suHkk1/QetJ
SsC/ngJORjOmShqAOtZIMo3mYqPOXTAQjdzOMDEKwl6M37Kj9ayywjEQUIR+Sn0+ciIY+typZ8YZ
89ByHBPjNLbJ43DDEQWTOuw2sPeP2uNfH7yaSJibo4ZcFHJWyeaBQ5XmhXXQMzJq6IWiBqycB/zG
msPBDr05MCBZ2XicJILDhxPTO01ab48n47ydk4juv75JiCLKorz5gJ0TCB4JVxQ2BIWRwht831Fv
YsZK+DzQin8AduLjFBNhdopyUk0oQlDqz0wmLXESFoRlNnZh8dbNftTGNgHnjgrhrSYAcgsTetZ2
4IWzbStLYTkOAwp+OrbxqfB/DB2EhjDZNe0G9rvcDqmszOeO2gH09ZvW2KcKQs0bc8D6JLooGiKK
7RlvDt7CMk7vC60s9QV1/kh3ti5x3Qo5sQ+Lrq8LjOO46J99SHymmOn8COEHJeA9h1wYvYuvDI/h
xvoSjYzjwqSxS52Y1+Qyum5iQKj5MPTgxeZCYFPZCxQhLGl+TrnksZOKkxobyLb6Bvlccknj6SXF
Hb4b0A3apHMarApr2P1vOZoPlOS4JR4nSycbyHp01WoHC61DXJ3aoThAlsUkwWV2h/K9UymZmvoZ
WHepjMMY3pMMfdhXEdkn+bdmhdX/Ti0O7cNGiukUvXnIZaePRTizYLQhCqcivaxW0AyGXblYE78i
aCvr7jHpBV4CySJ4zM5lAI4QtpyqR++nmpu0bTWQ5eRlaJ2h1aakInHo6es8yiZg/2Nh95hJPPIl
2BNbmKVQ/9Zi+IZdmy+W4HXQ6c+cer1PfR8piXop8qfw496HKHV74GkcAVrAEEJmN1Yxh28JzjRz
paaEzCW0tNZ95NnrwYv3QJYJ2K7U4pEc7dxbcOhAXV/7c1davCQBzV+kTIyZ3HG0mfsSvyVGLkxh
OytQ8osTShSzXUiMJqaXRdZIfd7mXh0ulaJMfOLCQbLkBIAxHDzgk2+uJsSwFncLEBMDjf9W3vIj
joaCiVWBu0IDvmKpJRgS2CLViycOja2bT1gMkk8GuVBaF29+ACi6p2PZRbJgT9BBlUB6JopbcyXn
kKLfFQncnY9hBDJKG7KmUO+ngJyHoMMxe2UjxIMrEgjecnMdKbbpUHdknIq+FTYGUOGzUmpiLM1S
5R6QC7+CGSkhPQ5cpfBi1GmRss7Fx59aBhbxBzFEQAdBxY6ZcKnots1v36+ITXV10s/eB/LXkJpS
TOuaZuQz1fcIUXvMowjkbbRFVOa4yqtGBnGx5C8IJklhBZIht37u33byDuFSkMfVpMr+0qV3/L97
W2LsuipTR/2cG5FhcKc6A62MaS6cTKIS1FZi4DVsL5B783EfdbAl/Bbpiy5Ei3pciO6zqq0zKHYf
4yBX/XjgPGsqc+bXK8iqn1FHr7h6J11zAAmTyF9cvcE6ZUtGPv1XlGracxZSiUVll+s/2iY2wxii
7FFutSQ9OgUVhJWKPXvhdKfdpJpbAuCmAUTRsgnD7FMTgQx7C4JHgBFDHotrBWgnOALclEWPqege
x2ldP3wY3kVhc9zGnKCIFJYDx9kpsfVSiiTUGkoPLqrwVG0OLsB2n0De8N+1quXQXLK1R8k4Vt+C
CxenXDWIDDzK93RXA31Wp6+4js05QEwLwCAKD3FQJVXFoms0pyhU79ASVkMFbg7eRIUK5jYIoc6q
4a/mzoiHSU9RlA4Y3hwv7Zs+tpDRNTP4G8jxllP4IuxcuRNe39KkEb1mssVT1oX/A0l22QfW4NRQ
DVUCtabNCqWaT6Iu0Qfp81J/b6fbE9m4l0WjlDWFgfYApHju0TPn/H2FW52qRp1wXKMF5hv9KQQB
VSZRMInE8kg5SZr93n913MLHQW2AKCwKo/ttm4j4fd2CfEewWSXYGPrgJNBx4U7nmW80tSzjpW7M
j21jGJQXi5cYpsVuG7HsxLGFfMll2UjXjvL/GFfRSQ3eRbRUGXqvjkfIJjSyYsE2WI6hrf1tjRjd
7Z4OOJ6SI3jgRbZS+rF6wl/dbMpDVX1qMceMZrpL/J7Er1xkcaIfhHAwBw7EY8LibUjhVKCbO2HZ
7DBrkR1PabiLhNJ9MvHmrwSVrVuPv0YUVVdUIzoVHVtQc6UH6ca1aEtGeLdyhAPcFOPvOmkTam0b
r0RrTKOewahhQen6G/ZtV9DaeCL+vMDtO07qw0OJtgFI4iVdyNEjI6tLiDR+M9e6y0rBn+A0GSQh
SidToAbE+7T+2dVcFWez1+aKUkmOZj90++iIkYaaIlMQz9Xwdec3gWNoaX0wAOTYax2GTEEQOTL3
3ax+Uokk+1AF2/VXuxu5OUX8W0EZ2A5UA6YtE/kRvHOUSKzuQB5OfvMhHTekKS+2JGXpHZDHzBb/
ZtR1uEWOY0JAnY4Za9gjk1sPGLsqhv2li8762sPhItR/IdUUhUh9qftuI4jMNAYsFJE8EDMGR5OH
c6NGqSbofG1KeB8nydFmd8dGOT1GNuH3mvQvj7k7Zp9Yak4rLagrgG2j4Axy+V/HvN6qn27F5EMU
zMdMsIgLzbD6Sh36f5Ir69gEzi66ydd3BxPSiROqmExYu95qwB+UqDfT8PxccyReU1PT4WCPajCN
X5mlHm84jtxCcmqLVzoYFVh1J7/RzpTNeP4qcwlSUky4r1rPFPo6s2knt6CkZ6qzAD94xjK0j5/O
X89k64PqvPg3XSL677JjDnZWlENEaz+0kjUfBUrW5hno65EmJ4ByW3866Do0wzGryJXWBzb6/jr4
8fDY3Rxt+GQPN1zBFxk5H6zRaqpIhGW/rf1bStNgiJBkzXCisdyuLrowiJXH+YwNqhyuhtBmjC/O
CgU/k7hZT69e68yuRLIopGN0fXLTnzDSv/x+d4yHO2urIbYMkvTq7MCagsA95fKq/ETqaLkgWmZA
d7NVe4m6MB8FrIyg39659PcFqnYFcr5QMI1ZvS0xMAFPMHtA8Auod2Qstfk6rjskYw/beema+S1M
j6znvXEBVChAgStBqZl0P1UCeWB4P9SK7uHUc9WM7RuCeLS2HtZymBcXZFk+G39I8fSpoDywLJ3H
Fhu5MjRy43HA3tlpndB8gYe+NHss3q7qBmAFnvrL3w9xil1bcOl07L/o9vRiDRn/wJQOaOAINvkD
tYUxHf5VKhh7EDlkYIj9Zw25fqK1WWsnwd+NTo+Xxe3VbPAhhPGTb4osLrUfERVvUJcN5wYOL+GH
cx/f/gDejLfxpfSz2cISP6Vmpg4dHObRM+2vkUosQcKp5mRLkFawcdD+GJR2/0xR7FqNbq8Y4E8W
72c9yFOdY8wUDzXbKKxeK4wktD6tGufGIwiv0+9lLRY03TL+F36UwgvUKnX/iPGR+3a+myJJMdys
uryHmvkp9+SkkcIxtFT6KySL5sL1zAOEKuVaVMUt5aabZMrx0AfSBpyN7l5e/BMcNgqgP9d92xhG
UwmcL/x6esyNj/72HMlhJlW2HugPdV5E7XDRxifrUvvXchxYBPKoCaC2EkzRk3vkGlXB041pTBtL
aUFd/wFUThoNyW5FYZmXhCR71MPmJeiZiyjo1k5k7xazM4RZXB4r4XmPvE0/ZSJCHz4eD/o4L6jH
XqcXuNU39lY4xIaR3Z71jt4q6uI8aMAYHBbZLL9/4vEYTAiwqXQJpJAg7qX2rl+nHIH/TI5x5YhQ
Qt8pZiaB2ZWHTbV+04DHc2DMEvBk4pB2b/jy3+nAg4c2LMti3BCcAfYPjO7KAH+BMJDL06U9Uq/x
CWywhsfeaandyN3Q2ygYxVwOo5+3wnls6gl10KrFEoeCcpaG/ssqCT3uOTzDN1umyLeyeiHFnEEN
/0YMx5shryJEe0gz4FoT5vs6/HlEOYpcRlfE5VQCL7bD+/2V27/M7OnrTc94U9b/E3Ozi0yRunJH
nKa64icCMEJnm2VK++0+lZi4J67s8TBGE6/Gl5KyiIjsZumg476qgDjOScuQ6lUZPdxhnjBUUFHJ
ZZlVURpbGrKAghyFPq0rbgfBWfbvmmmFEiQ9WuHPIC9Uzvty/9F9xvtDhmAYe7HTtd8OhZ1rQmFy
wGaC2JHuSV4EMYRhWqAiLUVlQhPEvqrDDrf0eyrpZVA2n5k4DjavbMKg4lusoBorC1fe9JysOYj1
+fXcHmsPnduGxXHpofIl1mb/9ogT1IFfIzqkXyBfvwsSVccDTPOCtclJf0Auda6H1tFgh3nd8zub
5+qge0nWKDWwRcgUJd0wSPcFq/x178RzMIusULFhHfloM3lBpTHysGDZjSUIRtHmMMJ8M/HZiTj4
Xrg0y7EVV0KY2gSvJf31V2aj4SWkM4znP6DZMfXVjrCyluxeGC/20lX0zMm4HDlKD5Dulqrsn/Ax
a3QmE0czjaRTyzQ2+P0MYapVMVEnInRwWK/94gk4jgT9gA5n1tb3PT3IuxRQlwOWnoiWFKmO+WUA
vgRM6FfY5Mzs9kCAcexSytXq4LfF8KTjUIFegIBQ8/C09rhCHj0IhafZY56R0gAWw5PuRsNAciF/
1INnWhDaNsYfsGrA5YJbupN90TW8FV7e+SRwXps9ZJYLOLagJg4JGzHO0NH7SqnjvOno0RH7ds2o
JeJ6APaZ3wcT3Dc5VPq9d6yF1Wh/Pt5AUI2EPvES7xipKDtxeSE043+sUV7PrKHKbzdUO6yZsjML
PgbFbx55s8PHuXmO53VUKMS7nH38vRzbVhgSnOmlOxEvtN4M2C+i5QKGKGjhJHXdPGZysK87QRv7
ntzy2nO0xVArPqN65tDmalK207bX/EZh/E+tv8MvCA47AVAgfX2BVrzomm1BiYfCYU9AU3EVo76h
4ANtxnFVeKN24FRMOKNJ1AjPmeLl4czzw+x5l12izGnPR5eW6P6X0FVuCOyQ44iiQntH7S/lOSsi
sgq9qM8xX/attE2QDlmZ4MLhzCc022Apb5GBCfyWX20RJrf0svKRCytnGvUJYyu0xFZ5Uu0h55wA
M5SmwqQ4WyPhe4iO56+7uUAdG+q106hexLIoOB9nilRV5Nl4BJHT5ksRTonxFIi3wEDDMnUhJroE
bPKkdpvibKe9ZvwSBRO92/8oAcnl7ewy/mJR4cN85kV0hIce2wnjI/L47PDd2Gomk/HnRCOaw6tr
/99h/2jWSajSf9i6coEfcDVYegUKkbRAbsKBXlUF/LZPrCPH8+zrMR9iCLtuQV8QGnU0BgkzEEqb
RBm8QVyI0tGHj/IT4ytBGNYp52d0WP0tonqSx5yAAi4ZaSHTf5J5cACM1Az3wE/voLwRU8r4pLJN
iqVCu7+8ZD6ZyOiqat9fsrYwtiwMItcyPKKX5efZVa0/j8UgsnzMXaBC19RNlLMHVXQFx43dLiKm
neNR+Iaqy1doCE8650PYi2y9UFmgcVwer3Zgo3ezZboE+tahxHz1+W8Hvt5y+hCBgySVJF3tf4fF
rWf6w07w0G69STme8FXioQ7xTviCpwDsmgfhoA+4ehYYbNJRUFJUwMkyDLTR7N9IUpulugovOgg8
XEsFQQKbtWIEityjeabvf91W1l3aT68uXa0JDdgtrizDKcbye1QXzQ7cQ7595q2LjEQFXbohbxDd
xIEk9A/LfBA/dYQJ1WAdxwAvLhmZ04kb+TRFLe6AjGtAY5q9BX4tY3YsM8a3Xj9oVqNKu088g3Ym
mKVOYHojDOeoGGNE2x2gh0WC+jzKurjcqnKS4XdeAp0ckXDBbliZa/dLzoLtIy19LR303QJxkmMN
AIm9jvhC8vWVg8YvwbEb2LYcUyjgVyPdaKozboeZ1ZgF/MBohyJihkEkEYRZbfQS+d0dUro8M08d
+BhMKaALPYgy7M6v2pnV1lBe6WJswm8o7wry5QwbuNBL5/vgkaIIFsqEcqJKDOMVVjoU2PyCGwjG
GI6ExjstBbeKnHG6NJZrJhNkICk8HKhTcaedZgO54EZ1LocdGkmV7/TMHIqKpYiNIF0anctFjXIW
1oXT1xwAf9ZXgQJlae6OUg9b344dxCtvYBaGk21zmVCcSLOsd2kXmd7xlvYeFK1M52Z1Sf0Ymvy4
LoxhdqBbjK2GbOlRw2dvmbfhmThEL5D3Ju0+cIIYQjXjADI3T7MlJ7KgiYz8T5xK8iXNZOqgcIHw
3bVzExDC54oxz7xzXE8PenHwMfBcn9mHEYh0AQ5N72JoQ7n2AZf+J71MiDy1XoSyu4h3p5wvZpWM
crMnapy2NckcQ6Ih7NKP4euEb8P7fBdWwLgeEJP30gk3bTcsno/Fi4pZwJkIbjdHjphHmiwdeccR
kiWh1zOcM19KsT2LDcb+ytD1x9d5RhcmyfozNinNwtNumJdX97gGntQiJ0l8Igw/qboJ+qCOccSi
g+Y8wDp15yitUmEefYMO0SEwfvyFMjuFXzu5Mbk3keINbKYRr+9Yh3hucqFEs+PVBa+Oq2qI4Sr+
wlaLlTR1PDJ6DLpIIaH7dRChvKfCooMjY8/sWbOTkhcbL1B7EVqesExx5+jErO8VzZdOvhTNfiFp
QcZklb0pmhq1C//LE/NuhNyUgoBLef/ihX+8j+s1kdJPm7SfEYnyXaSwOFtnBPtRZyiBrGBwDrar
YoQ0cAI6FKEoQNVSyFMbrOxDnSDgdicF/Zq7QppySdabrcGfWIbD0xII4gI1nW/vqAWlnfBuCdr5
md5T3IISchc8qRkbz6i+OR8Hvlfpkvb3hcr8UuI+4Jiek+rF96qDuDOewRoWVveVJ0LCQPQ4n7vK
XxmITLAxXVJcDS/4qZJLv2OyCbJ4M9YAIYlfzBghN4cY+sOpnsmBOxvPy3a5+za1e+kAR2O0x8K5
+QOFLKKXniy3oYaUnw2/3PBRui69rQ/XO1cTTqWji1dQT0SjDV7GGpsMnezaDWiRaIQUxyE4VHqk
aWwvEroZyBuMG/RWeEKFb4Kc7oJtZub6QyUXy9vE5aSw5hwEHL3jn4zOO3Eftc56lmAYPFug/PDK
jPRmmy5ogYCBZiYhdfZ+7Dz14ksNSItxUan5T/rQQSPSfcvtgQBDCXD3YsVdCJYHKN8XjdDay9V6
hX6LRMn6nzgM+AJMKNAlHSg4UA8WJNapxLGOpP3h89sUFW9FK9oQEKy5b29VJ4VAjeWTHP06DDLa
ZUlGu8moNJu9xCoZSyi2Avz0ek4L62RHEFVEapE11y/A1dNrYMlV4DK+rWKFKIr2v43bOHkkmjeB
76TT+G78oJfSZ6kXJSXohZLNWBb7dVG+p74vYiKt+h9JrzXYqjCcX0aFXaixJPnFsqzq47j62ps+
8LiZLIe8qKMeV+fNCRu5/v1HsLOeCwX2qGFQabDNHeZ4L44ayjOITXaCzUiS3z+XaulRL1MuVznK
3PhbmSOZJE3zZOUF0g7B5vbJNaHuyauNoZaIBMmhlJFOr/wGxWVMICWVRLN0k9DDizok6FJcvIA2
SNKAToGYYMNgSTT6RqmvSwPwTNPibhPFnIeVtrmWYVMADEvWkiWC34pmoT4pT6dWmcImyZhsYIdu
f3ZnCS6bc8CIJsT/Aobnd/ZNSSHoWhKAAk+r0gLNF/Lvd/H+/OnQh3cUqfHxiddwE4dIQ84fDfCh
qsRCVRCgAl+HXs5AukM0s1/vOegMIPBylodNRZttrVBZRRDtdKoJ9IGG8PVsVZTnc29N+t8CABhk
z8rx2fCn/6aE34Zsq1aKfEOK1d3Wwhk1TjGwoCgAlAoHoT4M2aTYBKHIOr8cjvdFC/AzOsZEeNVc
gqHjDiALc7g9DI1bPlG0xSikelE8Oh99mDa6sxg1SA7mOgI4l+D+ZGd6aQV3Tb+sRnLNoCeg/OBL
E6ACmsLDVnseQNh+NS0DK0oLnaFA7iOTD2h5K7j3fY7kYjIMfQ1UrT2RZLOaF1rulb7oAYEgqyl8
1dEhihP/ffJM5nJCtqF4vU4R+FYTKHZRfOH++Cu4E2wg5OXNkwgd5xMLhpgRJ/aj8b/wWfWTw/6R
oo1O9f1cSIDKcy09rti6OZ0zIAWYvUwDOiGUnUtfpZ/ok7XehjdQvEUhIk2DYUxc/bCSLMK2YRqO
4P1YDiDjzMzDXqyaublKpO5Ww21eq+jSnIA/GnQstkxbsVUXfiOApFEPtASp3gQnnQhYj6T1V64s
zk2eMj6uGbDy/K0G8UGwr4O7Trldurbw8+lALKD+3tnGj5ZDQy/iu/TXp7grRy+DGsqXT/buOfZV
0OUaxWJdqWKSXl7B28VeKk15cYcHAQFFrBJT2YzVEXc0xwy8cdhDbT6DAJLlzni9jHD/H+Ykn8dW
Z6nJwqg0aAGJ8poAQfEwBWXL+FF4kYHcm6u8poBuWSz/04Wfj2dFOfKWJaZjuPjYFpA/MrkUZqw3
YtB34JXMsxPLmNb3JvzWZtAxs0MgXaAVdMRy/phh41RWaPalr1CnDVzet+IM0ZqSwf1ZuLOaGlBD
eZi3A1kkGcu6S8gk84t7e2+UWcIbxnRSJINLAZQ53SOJEcCc/+kpeWlQJWMBkdtPjaUL8baGPP2l
XO9rLGOZ6DM+qYAazGnNRVlSQYq/d4VKwOJXSpBGiKTFSkC7n2xYsWWyrtKeqm13tXjz1UkqAU+z
D6Cmv61Ry2fWOCERLxmBjOm7h+Jbu1huv8eDZUMvTtezXviPiZgrxLJHpjW3hZoj4lu7cyJQxMnE
yZ1QEdd6TQ1qQ6Qth/tHsd3mtLlB4zfSqEgUvxZycoKdpWaVIPwTBhF4KNtXO4A2/dexw/ebK89y
IE0ue+jFEAFwqKnI666hgQW/AQ/FEaE+ZOxoX6AvOs5QU7k7cR5VtJYTiHZz4g13nb9Eh1M3JFT3
vJ3zI2A5UgAj4M9dYPsvtN1pP0kjwyFmtU1SaBDMRaPMVQ0gRIjwyUj/CqU22MCa9uz1IT6NrU3q
y/ZcKYPzVKkfelAp3ZLw6rr6WlL+ARV8QxcmkrqCdkZPS6Vi58rgs9BS87RirHIIK0VDdb/gnfpe
vvfGq/8r3+5o6qo4TkybwQowx9fHHDnuh08RjXHd1NEkL4iquEMLbANRqFcculEln3qQMDqcqU4d
BLSbX+fPezNSWs/ld6J4tjuCMVc66MZjoRSbAYhIBKoY1Y0ssnXEBaXdCc/XRu5e1bwrTgv3q0a1
btpHj/KATKRKB+IaFhl60NzgCKq8tAMF1Ue4/9LXjN0bdptKiRMJPhYliVgNmcUhLZYBwzW45k0w
vVqowwvfwtKGXpE2keIONnhSBRa+Vm3/13FcSC9msGEZNNgSlESr09d0a0q61e++7XKYq1Ov8Dc6
tMAGNr8Q+11bjXfQPF0kpJ4VzZHj6DM6DpdIT0k1KA78ibxuH6q4Wq0O4Sn9c0qgwnXDp3FUlgia
fNXD7sgCplT325MEMou+VVqkXr3X0ZmAPieyxY6fFmgHzgyChGDxiFWXsMU5OfVc/qlD8U5WTJVp
2DrYNA3E5E8ZiM3y2z6tR+Aqb8ziKKOzk7ItNFn5fnm5UItwFE+xoMzvuRxCHkQCLQEz/BoZ5xu4
zywxvvHanISy9L5fKlOrkSTq2N+cj2QIXpzL8kYR/P+2NS4nncKwpGQCZkiexi3ldk1qjgSk6fIG
ceAc9Zsvoqejr/+IZy9q6AUi4x1k8XFjAwyj2rktz+tG1iIAm11CtyBsUpYqZqO11a5yHx8EuF3o
kj1R45tE6QywbT9WwZpORfYlCYR9XYRJSgghxdte0tRrqk77NjDj3UYuUyROzUDJoVqWtd6cwx07
eOB0USgAo/1oSKfa22jGQddJCTiIvXqJB+Ie3dEUbpkitf0f5RLhcAJlGBzqrJ5+DtwzTyMc+0rf
iaXYgMbjsSiZzrmN7oM6ttLpsvnPFTF1VKsYCdnFPnHHxgdwKWy6cAqW2qkE/m+pLkN43pOiwrN8
yXJV2ma0wNXQeJLkJNcVkWMmgeMdJsSQHpUJKFG0XXd78m9n8qc1RC6OPuDzsQaHqT79xrGtYGHG
U90uKO5m4MTkCnfDwYUVOB4ENu8AqqbzZO+YHppOCGWIUUiTfMZd+TJyCDzz4GhiW/rXFmnkqxwD
vEKUMAvUr7lUHvuIv0zD2HKm4YfzIrYUxyFM1vPtAEH3i6gXI+6UAQ8HkYHvr05Btccjtu5/opTW
5fL2F5PoOqE+WMmwC8wpkSq69mqCy/WhiJTVfJRwWfsxHqWnHbisTS8hreZlBSFy4HxOmSi8PuDD
DW2GylJzY/hdnrcCDkWtJsVE628mjw0WCxArcloTnDFyyAjHtClPTzgCzv3E9X49wn7V4wWlEDLK
lJD8IMj5x6aB8SmXtTaPLQG4GP4u1sQYb4pi7BPCqaBLCQ4y3T9JRK+gGeAQiMfPEo60/NRmjoKF
mEXq0Ss2TGGPIYBiE5yTfsVptU8PnxCOAssbpoAlu/uaqQWDSKRfLpIa118jMWFX/4uKa+Q+8KpZ
VU5HvhpX93/yC6lQn85FYHCtjWkKuOsnr+THCZoS2IOl/UgfAI9J5Wdrk39XezbWQVFoFvsgpJ98
kRa2p426IpO6S5CvgX2msgobVE3NUzZ8UVBlN8edJyR5/b0Ff98XhrDoj9LYjeVbScK5Fxccjc4B
HDFXc1IwJtypXg44oxis22/z6xBFG2DN2OjdCahAWfMD5XAo3jXPL6RHBseEOpNKQb3sMvjdxULa
E/+ha3OUZD7oBzvThsLYR9W7147zU5rkF6k6YZlMu5spEOc0t6mjXoxYyKriMo7MCP2AEBWFv9CJ
L72MLrBHM8+3bzyQgQL4PugEJ6oRKuAevGy8dqwQJRWnUQlQ3TbvFpgggdsxqQYZxjegN6eiMJkV
45RoFTFUuT0K483974DGiceSC+Rta+5rh+ZMyqWeM+Q99wiDxY1Im8DXCNhAFAPm/SP4QzkGwR42
vF+8pipdOfRbLqaC+KIJsDW48niegAOvKGpmrI+FjtVG4O55drXd+Hxkzhm5d/TTKXJDMfDj7lX+
6Cj9I6stImWQhD01UaLDn7bdvD+rvUI48KziIodoHBhxhUkt9vzBczEfP4LuOPuGr26N3nYx0aLX
Wc7/ZP+BiBEEV6zqVDG1No3CIhKc3MPzy3/RQkYKSHTolT5byRsNYQuECgCqOtS4HB2Q31B/8Lwr
Uaku4tK04qxXeh3OLjq59hP9OBQA5nxUEXje9LcNfk3+47aN6ORD5h3oVxYPKw+dF9RL9WWlqss3
fjKFUSGUhNUNd5RsumqqmX99htvBdXlKQ1AhvU1Xzl2fVgCludbwjNVuFSZdCOVWixPfEhRp1R9W
9pwOeUMkeSUZs+EU2vD7PEjx73lhXj1J9JTQ0+naoTRWccYaqFwh2zDRjiFUPATv4RCxHbtjJ/kJ
B+QNT7Tk0XhkFxsopqZQKLuqbbkmh3+a85c0FLcw3H0lhKLrzAupMYO9NYTnqXRti7gwfckKd88J
nKJQQCIgAG+Uin27f65fFYaMmhpti+bKxQZ343vWLzRhg9CA1ZvpHIoUT4/1URzFl+vWTgy4/l4d
reFAT7Ugt58WuekNbQ76um2R1PV8/b1KghqyVOSSnCZsEklZ5dO2CI6J5dCj1D6fJBOgCfv7hDeT
gZGPby5h/4Vu4+5dk9goh4MVV9Q5d9wZRUIAdTQRkx0xKK0ZD+8wVV/rDB0FpLwUOI4ddxhOWbpw
bY4j3Cr3GainLoRj2X7NqM5y1qhup50C1+6W2SexmVBY3G35LkIoo5QBOicpkMEFyvnrGePwXlw1
DHIaJIOmUihazmJKUpQIK7qPS6NoIds7t2PkVBNMqzlqiVViXyyuM+8qrZlq9q7ZX9Trc+MBl1Sn
Ir2Jtesfi9YeKduSAJJs02touEOAf9BdYpSK/zGKgdlOo3Ex9m6NUeWrNn7XQSc2sd7c9BRR8sX+
2I4gC6MB7PE+D/anEF9UGL3v6yzyaZioT2CbrH374/K1Jjvw3Vmhox5OS54Vn0RJt2QwGMmVsBvK
LFdfTQiUtPM9FHiLIvCMyRyJc/wfEPliD/6tiQ5Dz6jUGQDDRlFQJxuSwK2bNTXCyOwY0qELdNlS
xtJ63P+4iWl7h3GCjGNY+bYdO4d+OjgBL3U6JzJJdJQveE2Eo/xmT8DsCfspRoujzNCnAto8p76o
EIVjIXL4KevRw3vSevJIDYsPMMrofvWss6//LQHFtcDntB3DIfDd9C95vscU5pauhKurgUNK3Rp6
s5ydmst7TAZgZwrnGJErVOy7Pg+g+vsrS5kMv936ChLMujuebRRareu+J4TysZ0NYJ9nZxlMOs3B
COmXQXaB6skASgCACUGp2m0uag3aA2jbgbLeFfBysRXn9S7CGzOQVIzSYZd/mPZgrhSJJDVyLDpA
sI12wcWyjbBzu/xN36P3V7Cc+OYizyqnLtkqOV6QpgCAWtbVwvdJDcesfbVeqh8E/ZqsqggZcr1m
rmEt2Ai31Uxr24ztaQbFb/sa7fBuH8nl5mjO5hArPDa7w3ZJHA2yAqT5yk7bX5b3RNgqRBeAcPwZ
kerCW7OcPp4JOhK8mhpjLDCg6iolc+ic5ETlscPDHqpvyFKb6ZW6+/sSEnARG6/mfnywLu8Q6OyV
USxpH18U0KM+T0Kc7GOeGQn80aNtMOwJEkRpHs5gAVb4asPXQG39MGl1ANeHw+GO2Jul2Wo9wVpf
3ytRx56sjkiFAlDistE8k+eFJpCw6CGsW4wONOFyeijRmNfD12UuIUEf1mEFouUe36xEfHpdhdJu
M5Bv2gQ08OrNrUnV89h/in3nA9BQrwHbHxf7z8/FZJDbqVUc3BPZHKcX9mmX3H7zbzTJQR3Ntzi5
OJEUfwKKTnd00+xK5c8wSUxTf2BoJvEUwTHMqY9hXvMCp6CPwwl4wgJ4MNl8EbldbR5J0+80EC7u
dDwuJ7HMqG7a0LoB6EmkWnv40f0R6HaUAdeSfUZ21TRsUDgbqV7H1k9t7zP7vqJ64NUdebJ2A61t
rRdJSEJ1UcTbbhhiHLhyVfGrUJFxm47Vgk1OeWShNlmGLFwF6vlypfxS7FPfSexzn6uX13f3Mf7q
d4s4TszC19KOXBnODlnhBQVINptfEv3GtvwSITaCnm0dqgHVkveKr36s+Z3aOrq37eVgAkLtWBC1
LZBDtot1M7Qu9qZ0uV4zDZ4UJFa/E+izUiK9tE64rvEiKaSjf03ZkqEInzobKZMygKwKA0+xpqlQ
xXa7b+dimcAoWZVFgxvwDZO4fXIjslt45ZiY9ZJwBneNESTdP4/GS0de585bmJyqrTXNbMtETBPr
oQcZ+vGBzYhTGA6zKPD08XiH8E9PQDM588qaFZWPTznyLTGSPecK31+9RXKxx/YStzYrjS6v+5M8
ZjruQBzT4OenN6WxGF1PMliZp6o4dxMjsWZ59ANbLDmhZNPLdXAggpPrehGD9s3Yp8MQTGn3ezKS
eUeBcjk8YvCvKPV52ehWk1Cjw4WJ0PLDG4RRmiFPLhNC8dwGDScnfEJ62yZvhcQGb+jfsm8UYFTi
q0V9srWA0jSzfEmJhmFc0axfDh4hJPmrdUnbJQujuxWQfxUU2uGrKRr2eR4aPzKfisrRnDZ2XyJC
sJMdRZhIXiyWoIv+3E4FLLleO/TEqbhW+Xhdv19ZDL7pvxsE95cLaOaPM8NW8QACYnoOrPrP8i7x
xUPh9yGVXe9X10ZmOXTUOUPOhtiooM4s3ZGQmeLYIyDE86xa5Ox6KlCJN2Xg1I4D+JTPvDJn2eVc
L8JzBuhijsfmwsMogoUbuv1Q2V8NuKDX/7ZDC+ueN3E1Se6yt/4SYWpZPOgEDhfdrOFFsawYwIGr
V3KoSUmk4aby8sqXN4jPI1+LL5hOZs+WHjR9RElxkJdeB0OWGySGSyAN3Y+rSshMQE7Ym4AxT3mY
cFB5lYqxvs118h7ZM5yQNEt6mcdgO4TvCW4g+6pHGgTe7EfisABZ1ajvsrh35idk9coFNuxFYOYb
VCMJVwuovyXyWeLwfvHsH3K4IbhlifQETRAN40zd+LN5SskPjp9l2wWvfhtmSuXCpF5Rvm7FrHRD
DDXamC9FwXYqRTB4tQ/UZhPAeU2Obng40Ljr4cbCsPXDAsI9cN7BGpFacV4dhhivG34aRZGXf9Dw
VdN9kxVLiEWG/Vx14fd2JFCdlpi4BCj5BVhfa84rJaOUOV6ML3l7xK5advNbHUXNcifb349/eme9
d2U3EXa5+fGuCWYgephSSeUQebDeJ7uMapOOtU5m8VAwd2/0DIVRbzk21zx20j5FopgTxUhnNzxS
JnC8xvIezzn9qA1IGNf2QBMLAnZgEESA6vaz35kvmFrPPRgZxo7EDAd9OqWhxqsr/u0lS8+ZIxsq
5I/ueR84OT3iS7chu1astdmeu8s+SmwyDBS0wmcOdCAn4L958xhzBeNHKVSaB997gjTzfv5JIehi
0OlAvxmEOUQXpUZuEhw5Xzklf/Vqw1v6AwnKFrWHQsy65BKtV08E5hsXRYmcsxzEEAEHCAMs2IYV
Sr5blgVS+oVpPhaUV/32vLlAB41zx48DkMj6mgx2fF4ddAnSKfn69y6GZc7BM+Nj24AxDnkiW8Rm
YpyZDYd2KhY7IZjt8iUbIkk2SG/JdA5IkeQqgkC1LUWOTFtWJtOd+NuJxgDD6DUNJBzzSPS/38PE
Nn9ZW66Jb40kivsPuRmK8hNXD9ncc7CSaDiMYfQXsgr0aUwPzbiQCzIPUEl+OGcVdI1qKB8y7mMY
wM1rwvxfiWDZeD4k3Ro4++C/qFQFWpLuYyHNND2abWJGXBDXew3NCixjur+il0rk8qD+g8/Gx4We
aBZemvpwl+pH5UwwUBPmidZS4QrGkVpJr9tJpDTBlenNOg7H37SKg8+kp+9TYwYax6JOCvtoe9eR
CRMEHC+XgcxeInUhNlWJ4ICCneTXu0J+SYfEWgx7WJ0cOSsOpeAzlpjWGawaQ+mSPe+/BxaX1hV3
2iXkiDWJRN4geKVhJzdPjeK/C2K76PTLLvR9iK9ltcV/IMrxSmg1ZzGh/k7kjx6iXD/2gg9lBIv7
jYuAq+NDMGvkQ3/frudBw3NQENY/upahbJfepuHUeLzdXKKXTsVTaPqAYYlj0nrjci97JM33y5Xq
AKQPagqU5OLcrRLgit5xo3cqTDFKR5NyY5SL37cORlGy4gh4B2++RMC1wX2wfrwkcRh5KhZo7OFe
z1c9u4GFPvg/2EZsNkv62jmhn50FuaBrVkcQlovTyW5VXlqAraBfR0thsCUHmVbNJo2KHLbY8NYE
tCuEzyw2lhWvOhYAnlvv1luSonElkl7fiGb8uyiJ3NLroTG2iM2EUeyiwzqHi09zmtZBnrjTh5Sx
RlshPDsgZHw0ZT0lBIJau+N/lf81qnYwIrjdf7X5Qq9H9EKlX95nUdkmfWTIJYBaILvbaq1N5jON
TeHOme1+de+rZS0WbZdZAaBAvU606l3XPkDctr+ecEBMtqIAO2ijyYiD/xd52irGw6lghwZCPtW0
Ej702x8xLYBaOkzt7xZ/KKnBEJrmM4nuwdZYugEgDs+LvHxqcQ/LTtHO3xWyia1JYcFEFfeYOjTN
GxUPRfvnHmYvh6Dym3tFulgsw2qd1MaocgRxijBX61UwxaNLigGXe3wxHDhhjFC3qZhZragbWdlN
wBmdwhRLlEnQk69qu7OBzu6hMNt6VwwN/+pitngqx5/mY62ZiI5c7sPyrsV3Kum7wlB5tDipxQNb
4PzjQegdh4nG55rIBz2y4sReP4RzjeLDTV0C467Lc+g7RW87T+tQSPL9Hp2rz8OjSNMk/pQcGLWb
2GVIECiDddHAxhmxNM1rEv5EGytgIBEBG46FTQQRxNWp+Fwb1s9ZIjnkP3+Y0FZYUhUPwvjRwB9Y
4h3YJSmCWk0QzwW0ud3mFErDjEww8FPZGeRpVOgRMprkky7T2MhflGPCUq+SMQlYBGFy6AEx+zfN
vebegBBIKOvTnTtPLkMddbNptu8wFqPWGLYiicQbnBFbNKSbpbsF5aPnetJr71E5wQG4qcnWn4ZD
2Kh9IXnx+0gRdo3EsrOSb8aosvv5EGN6v//uVztfZKLXUGBBX3UttOXHvvEUD+BUUkl7E1/FYq4E
PcQNFnk1b/EJRSkCSMAEeePjLK66J950Irjj4Q/Olk2X2yNQYsBnnewGMdeLB+T0UyxJAKSZFh6n
B+ALBrWmxFLIA3+p2YzHGdPBkBZwmsuDM3jEiHD+wIngjFrnNHYcRAMzzmGzXMuMlm5zjVEEZpQe
jeWB30mv2BdNXa+dCGyn+yfqoO1IEI3aPJ/AdcXvoOJ4II4wKhh1j/hXckiT86Hc447rxwoYxIYe
AaPgOdxe0YEi2FhIwZCurUVYH51twDcjej5lktJgLhiJX//0tENc9SvN1Dacq00eLb9zi2NTIiqM
8d0CmnaM9lR/vEl3wTWrq37Y4lahlcpehkgvpIUZTdvrYOr0qZ2PXYdZuifqihcw7qgRjFyMJgqH
k5reu3kM2MNdPvUrAB1PJMsK5yGe0pRlKD6NBG0r474tbMS912DIofsDk9fzPXQAw6Jy3nhlvnRn
NZ9nNG+fp+/3QePePcmi/r9lFepXjck8oRhnWT41luBlDK6PEmGLi4RmAjpijfe9zcPww/1Wsvmn
Pdc7C9sNPZkekMgxv5V2P0QJ5GigxW9ByoNs91Z82Kj+Cv+zYGyYi0I7ds6ZmtAwmj2uj9dfBXLc
Ci7sGeTGJLnDjRA+jHptdn6rIsPfrkY3YaB0PFbXpxXinPb5lkyQ03aFFuesoRDby/1aT1VUkJiQ
Aho7kaUJ/p3hYt6dUpflAlkIyVYNsIvcwWDKARP7W5iLOR7MaFtXp+qYxZASGZV0XKw1rgBip+S+
8x69ynGApZyejIQofSQ0qjpEdoZec4/5Z/0qwKo8l6qPsbU2cnktcyMqO+ocwG2EjU9025WJYX1N
ILIUXk99tgdekXoMwzw2WB/RwT4RVa17HyhC9mz2swj6WblVo480ZpaU+aC/vocnvqNixdNBCU0n
jw0tCS1h5GwdIrrwAYPhFUaDCJ3FN0BgZQGEbkqQegEe7qqX0a5B2/rAyyYf6ab3GceunvtRYNLT
kRvHJK5V/MeLhZTh4p9T0PYcxgzEin4taPgNzY/6ZoNVUuSi9usSVCXaeQufXQlCvyb5qwVam/Ph
ZMcCI1YDObAJNFjlX7LtUuDgf5qwkO/+UYgNyNuO+whdSfbYFbweDqn4W1g9iTFPhUez63zk8c7B
hWQw7edJ06bW2tP3DhgkHJFK/SphcVOQ5TStR0+NgZpIv6lrSOEdw1MXzjO1BAntaGF4BDmyptNE
nkRGj5crcvdAzxld7ge7bVr8KYiGKq1Ql9HjKU6Fvgzl3Z21Py0ZGCdvIaQeNQKJBuJwjB2Xu3cX
wpSQ4Nd5gkfC0LvdzbkmwgRuzD3exDvcovSMUUoHU3EGXwLjDMJAK3wfaawwrlAPkJv1HIgferJi
5qCjYwD5Jp5BiaVqf0xTYRHlp1Exj2O89ZAjIqIxT1zlaQtpAh7RnBF0jrGf3Y1EKE5MMubTxOtH
1sEke/fG9kp+r+uPbpoA7mjTwUH3x3pv0Usk4HWnwowLvRst4+zRIIeRvynPTyJfiJjoh0tNspaW
AoFBUcLYKmky2ostB0kjB4h/EZbMMg2VFmekTsGxVNcxXBBuP1YMZZ3Xn+ien9D1vrq8uhq7JYI6
OQrZVO0OgStfamD2Mc7ruS0ekAplBWAUrWRr2BbEqL1QKSl0XtHEReXaGJHOzjfUWng+U2SKpVdH
QCTo8sR8dGqhwRa9nk1i8R52WYrtD0VZbzG1t1FGYR5Q+zo/rMZ5UfyPRz//jgTFT7Z8NkD3v+Vx
olzzY55z8HO7fkqT41Kz92P1trUpnhL1fSTWPS3ccWY+XGQ8g5LJV6SIQuU4+Mz6+pa1kaSpIjBc
TkRkm/ATe+523SooBSLQFaqMhzocqmnaHmJloBEDlPbRHFj+ClwO3LcaiQF4hCNcBQFxN3alG8wo
7x0fZGOfCXZFI1bdkqMbQF3iBwT/HycZeFdjwxKCpmT27Nc/XvT0w6r8umgAmjvoD6EN1o2vdrr4
to5YgrKFVLKcecrkPephQZ+hc7YZsksbN0IR5ApvplUDjJrUyzUI0wwmaFH/IBpo7YAuIMldeiiY
b6qd23hTtcKbamaibkrDSuqQOO47x2iMFukiYT/k6kfr8+ulBP7bPQ8OnjTZSsPgPRDeEJSBosAE
woUN/t4xHNYe2L+28C2z29YhogqVP1XPIPz2sLWA0gSb5OHsrHdvHsD53JSI6YtQgKG7hhKDEN3q
IcTxsUe1lFKChVydIx0gL7YP4DJO8UbBcPnZa5AZDkOoAZibfUSFVNUOKZP8Pxku53czh0Shu5BQ
3K9USAYzX76APken83K5um2sBo+NBv6yNdtT9QbDPW4LIvugN0dbFYJG5yX7RHB4XXS4NvKdJ7W/
B8D4886qblwXcW0HjjKkWk9O4Qrt8OJ8B8uVtggQKEMsNw3fdJYF2V93fb5uQ1CuDRnfCNX5/D+T
MhxrsNjuOgBjBW3DdvtjTWG1tDFlY2CRpu1LAz4JtE5eb9Nqvwy0cdN9aSNXxV4FIjd4+0rEV4so
XunP1PsxruQcf/WPvnRwBCOavRC0UlpU8rPNNraJNglKVhTRscvd9cdWb0HZfOWRxO3sEXDdfCNS
FHrLs7VArz9m6OE2/vTLv2jTza9IvVHJl8m0uZlcuYEeoNJ+8WsHAPmCbJRn8wzFIeSd1tclpqnZ
nz9shqkRoX13xFRVJAYMCC/NJ1IOzSqtaxDsHfROfpwDWURhokiT6FatuHQq28gxyqcox/S12n62
gH+RFxviGBvsK1+BHPoLAqn50tVexE89uVJdPYsQDWGnoF5/rL182aBZ8cvP0mf1kwUE6AVcqfDY
hPFUH1wsfQB5iZEOHJcdYjdoQzxkhxebbkd/+INue4EzmOftj/JXXriR0OdffmwK/6LS8bDCfBM3
TWzTVmKONy68J/oKY6Gp02AokJZWFBLkJiCpb8Qx4E6NjvbjGAMV3ZN0h5BkjrfxhPtCbYOmc4w5
pcFcEGZ3VPeTptvhv/PaiTWV7A6G8JwHSTp/IRBcrCeTjaipp/pfB5igt+XtRNgqaSnY+6QunKAr
f60ZiXT3JEnkcTFjodO/muSsln70j2gcnsZp/n4BPS5H5O5fdO1JEE4/lwzCCNrqx9Kk0LBDoTJt
UlabiPMN81tYnNw9NkLfEde6iGom39OKd/eLaeTZtdVZncv2HWbfarASTv9TrzULdgU5keuZ2n/g
M6RkMdy0M4a/4BkNJ5+5tcZDqh9Z/oWigJyu7QTQq/l9CYS3XYhnTT4nmbI8qsY41Ja5WqcjREYZ
Qph4eWvXOWXp662h6uUUXEbkpgkRq26qm5lVNqHBJD/jle5nb23Fy/5yTiYcZzWy3dPA+Mo6FsAr
nOOq9D18aJZR+AKWG1UqJZjO3Q6Zz84y3kRADB7K6wcD5nv3g9Pz+PPmGoJXBau/T5wXttMfl7GC
Xp4jn0HFNpUDNwdoacTYP9XThjXm5Y7TCkkbFUFzF7Ft/06OvxTPyNEsq81ZIokEzKY0TBaux0VJ
DDOzhL4vNYBrvo1GgwpjOpvcq86j1UG7cy43/Wz210sYAUZkbGkAc1Y5AfkQfr3ceRC5+hTNy9IZ
KHPaSOViauRPVCIZc8RpaUtEBBM/vR55CxRLuitNGkKdXDZnUFV6PvTZe1HjA+vc8VoTersDKzzt
wmmZL3qgLS79g7OMeuSxVY9Lcdgf9gMmscqzvvxiLgJlEXD4HDvjlUn9nRAf+xJe0zcGiWDH+eL0
AZTegk0/6fcJkeieT88YkM4WceVxmITCgi/L8t9tUdplrqq0Cucxn+nyyv2M/TEZkGN7i/BpJUzV
YagwBpN8wviot+FegutmlBMJASHRqEIdS2loLVXIgIIyEtzBQp61F7I31z3YjOuuUxuQezj8oj52
+xtMGZwdpU7bRQFpZjbHXbZqG9L/ySg4gAVMW5AAM05XCnStcMHSGYvDESSmIgkEkPY29pXUSlKC
bDIboRgnNGr8upo8YdA7TY5Uv4LIknyVhMAFQSa5d5nGx1NQexUN+4wqDY7QxbmcAY3gwDD1mRed
+isq/JdnNEsCowNbdQnQDESCQm82GTp7PjBb3wikptLRgydkEzSkdYqkuFUfFas3//a/41HZVUWH
tAknyuDa/cx7q6CW0xCPWm2vk6F80P9jmHrDVhDBwuuYJDj6ssnOHIXoD6TMFg/kC0HRrMWtWAOu
xgygSGmSFNgx8TaCTcMOhuf60wHfDxr+dX863StsPplg95Vm4XMImvtMah6hkDoGgK8tr+ZeZtP1
qfdShTDLF0FGwUQi86pWgf/pONrA9ZdrWT0dQOq31tdbT7J01YJ364DOvVwH2VuIOqGuAYWqpw5J
/fPHU8QxxMlk788wx6z0hDC8jaPk8G6pYLU/kU6o3DUait4ELWdHvy+YUnhTszm/kEEszhIPbIwF
zoecPX4AcyDvcV0Yusw+qjWNpiBSFoqEr0RzOH6n1pjl2dEqAOGIQVpQzS83Z2jtZhLHjlDodVHe
RwW3z+CJwD4OTW11mY3khENuXSF2xsjZUSqtr74iHHZE4Kyf3VocHyuyAAg3j1trtoRUjqVpzBPg
wctH5w0EYW3Pf9p99ZIS08NMgOkgXHX7QDrM6HE3dHd1iFBWRhVGtX9B69ZHGBvRx+JhspV678ef
LJj+Mj0OEY2zqJStgKBkce4e3WQXGeLJJnrON238YJzlRpWV24TI5h4vHhLU0EReAWHpZKHIyur4
EkNGjP4aPsCHtXwl4ukyJatUVXrsmq2ahe3YYezv/b7Uv3AnX7qRgJBBzw/Vn80Ox/XyspDzFVQc
pGuRblyIFDLrBt32VFglPJ6Lp1nNhnjZLzfFqcf/P8qcM1nuU597BJuFEWK/xw4t9Q3fthrBUdC8
6Kb2zfGrExrk7CCeuAVmM/IVLW4NSxC/F6IHxUEm5aEp1EP31DEKghaEN47x+CAW6fBZNLVTBf6/
5XHCw5U4sAWET1mX6AW+3HJ02Qed9/t1w3bGpVUAygiq4pdMbvFYPde7q33PQcfXG+bWI/KFSpet
ua648siPsXSBiVq6W2oOO3/FFdSxjPrCY5zCksTKX67sKMsK9jEHv5fqrqNaLdI31rFhCwyKfJ0P
1a+Kgj+yJzRcPYZOiEMF3p+Qy8od7FqvxmQYCv2ilL2FaeDV0y+hHu1PUem+X+SVD7MI+ZS5TVXw
xf+qf47WhAaFeSpi/GkqFinch+vii9Ba1w5pGrb7upan+g97NuJqTMQb+mowaG11MNNx71c4JUxm
ALNhu7QX4IGJku2+ONRD4Ax4tSeiHFIvejHqvCUfJUbK5l3FUGICniE1Ez1qpFCsBumuj1QTr/iO
OrRoYR/lej8SbRHbA3UwLwJgGVuG0+oQ0+gVn9D5MzJhGqnUPkEhKaUWtd6WWbP//R2aQzCcsgKF
JogqwxFK3oXUyStnEJydEzr9+wN0pG4aPYU3cUHmOr/DRSwj8qcTklocHu92nNRH3xkVbcxFQLEL
/tRZXyb8ACSjO+JSAzssr/jqFnFSQ2bOWwYLS622DeRO5P636wiY7MZRlzo6ET7ZPrQJ699RB6eS
qN98n5Q+mc0FhQ1SbEFlFCnglxxCD3S4+BkCjrISHTLIjryaAX8CExiskPoRTb/3P6n5QjC2U3Vk
loXb9f+95dq62/KORsObZHexx9nW4DDKD0PrngPwS7mTCrTKFoY0KZGfSzfqyQ8ykwsjTzxI42z+
SY9N2nunk583WMe1MllcWB+JPFCH/eqTyzEYmAq9gbKXXvvWSKlFVSL68B4zsVLusVu6enmPJSDI
6qPkmBeJhv0NEEItlEZUQHIrgoaHmd+g7ZP+kUre4IFM6ke68ntqskEYw3MkKQk30ohzz8WOH+29
i1gMEVGkAdMFabwYJFEj04hONO10h9LS7eQOcGYvHZyRfHI16UYzeLnyTuN/CPXL7z7Nxeq4+Ipm
wXnCwpZt5tpiCVSP3xPa97C46PZ+lVvHxrHOBVEOJncmpeVW46NCE5WhIYBKJMMgwny+YKxK2Uka
5vQZC6vsQVdaS9+f29EnO7xw+bU0SVlmKHUNDN39qhjcALeux7TNWXsUGdMAPTBtfDSZDAxhDZvZ
OmvCOGiUV3608YRTXj/OvsQoUiNZ3WeWXn2yRBbwxttRC4O3Amb4yVpHs37f858P71zZxSoJzlj8
IW4vFBMJjMRqF1yP+Ez1sIzvBfZSaEfa/kV2wbpB2U1RKc8v4skQHFqBMmKzYXfNbMRl2cn4cv++
Rsk1BwEU+A8X+Eh6fxvj54HdCmxGXWIC7JAVnnygLbOFW7dP3FLaj0wnj6jMqCb6rB7AxGL0X7xd
wu5mUCYyKEVd06avN3SbbTXvcMYzSWkwPVXws0xm9GeGci+2NfhdXLMtSLWfUV7YNhHTH3fdkcC/
IGsEZsM/TALflJVaSDNxtRmDJwWuAtI8R9rHK5gJBiSusb4WZoX2u2ykQRWiGRdIKWybn9PMdeNb
rVtDLBtYV0xF/uhvjdMkiVWJnoaBxU61AlBCbXMTmPUedBOaUF+nRlf0Zkv+yuYnAPJ+sySpk3C+
q94qXQ4aPZ107P62RsUGGtln3SHdpM+GCStY9KaBBviBz+uPX52/N9Jx/k46Tk6QFsXWeoiOn99g
WnC82I/HGZqiUvlaTtIsihLPwRsP4wauwsGHocxosuHLr1lR98xzlgV2IEIChDpwAxYYZbBf4QLx
N6s7TKA6LhWWixDl7GtCdO0WFRfdQjMKH27vigRLWGMYoZByRIAH3bqMltDJNOdQvgwfdlpmEuaO
rEAjaMh6h8b+GGOPC/19Znu89aYEXpbXNVat0as8coUbeRpKjPM0EXc/kA/vMDV+oxHiMi70gZJb
fsN5upjFKoUfpeaCjHid2dhN/L3XZHbEqldTbFFqyhkHDZyApPScOicLgcqqru8aH2gN9JnjVV5i
XjNCugZV/MZur8s8pxfA1wCEiyrtpc5nAaIGco7kBYsoc4DNxzLlxK2rpFMnGbnYGfmQBPC7goWJ
dQVzUkEqT3dx58rs1T7mUfgaIuw+ILdOa5N3CIN2rQbGFQ6AWMpGdbE2j9Baim/yg8YUrwxLqL1+
vhslDf5kgfE/qt13A1zKMKcIjxZZ0phFWuPiaExKzqWyUgHhnaUtYO9/2vp0oLeXv4pHKASAg7in
9UBTI4nTrFS+nC/RlrfqJs0gzolTXsir831JdDgqy7d+AAP6T8rpQbZ6nPRKjLlcWeXNaPaPEkcy
uxlKaSPIAZ3FvxXrgARCIdLwG+Qroq0qvA+Kl9oeHUko7n8SPUgyGXVQqwAYnQV3W+cUSB4wuHFO
b88jLQm1p8hzLbP3ypFVRriR/df1WWidjqdn2XcX2kz7Zcl/RaTo/H0q488NDbi1mcaYx7Rs3lHO
xXZK+jwz2OwbPjy5DFSterXpUOL4o/cbmyBr0YUByvNd3mEt0ZUuBKL00KEy4GMVJhV6+CbA/xWn
Buj3dF/n0dhHB3VwAcIL5N4gtOxV5EZlYiRGWfp6ThGTOeBEZZ5kQXmn1pOsbtskljcTSm5lTser
wNZJLSJKWXtv3y8PA1gIQNxGENMQzPf0IQHEQBMaQercBZY7ZelgyKIpoB+Pi4TsxUgl1ApZUREB
rqF/5v1jmHj9NQaZH005guOWagkDneaZesdxnyiCOHzFZMBlWqS5ODIn1sCcDjZXH1F//AOnVZ26
dmYRrYomkx0eExMFd3VxYwehWfZnnYZnl1hGZnbRAehmNIr84PDWtbUjM7dE9z2oB8+Szh7UjuWz
JYd2mVKXPaYvaoXDgVksu0zcMKQgahOn27FPSe74WzV/5w/efn9OmtT4h6BoBVVH37e5AoR21TYU
6MZfF+7VZYDAhVrTBTch7V9PekEyQtsR7U9bG9s4HY1VIJK1vsihsMC3UpMzvTDIXVs7Elcj5vxr
E+b/UnQKqUdDSv0mKhzOWvMrClxahKRLb3WSUVR+YBz+pVKdaBN08PZRkD1LDugWEuQrT0OexDvv
6OKf+OCtQoUoA/D4fB3DkEc5e2jeTNJ4C59HSsizQtyoeWSACSwnN/hvEmW2fwMQEtBbAsHKiJcK
IUdGPoVZhtLleeN77IwQGoGOVJObnNk7W1D+Q+8eoOCCSDW7OkGy76X4Jr1i+kESiJp1iYHwAWVT
MKFuOIh9qQDjPMxLQl984iNlzWqjwued56VCtPaxYHieoQgjOW5byrpMsT/mSR9jS0EmMvHzg8j3
wPLXzz4oWK2+z1mDq8LVx/91GNhZtfifVEECZbq1hjm4bG3FPtuGEVHJYBCNefGrXwjHKmPKXlw2
EdiuvAyXg2YKXxuCKQp5G5JT8GW/qASL4/03a8gMkrmauf+Qv+RVCqPHgovJ5QeiO7Zqr89wXMJ+
l6UIhS/+e2isuz4KoBQGEtmdcga0ULb6JGHfzDNQEkJQMTqL08O6TkoK0s6hYtF6usgJgCH+ZGz3
Bopwlqd9uLJ5lSHi2BqZt3TGwpVVpRh4EhGboADN1bSvZzYkjGb9Ht58yo5Yq/voaCQ1cSVrD7dw
WO7bY9JAMrhoecJjEIEf75Kyo0mLnS3MZ8Y/8mQKVycnHYB+VAzKUOHM5DqoWXeyZWVxW8n8sB2n
4+uxyYnws8M/pB69sLERSyQEot9InkVuQoCK6acqKT7ILCJDgf1znoJQEFowP2zqDHTAga17s5Gb
VGdNhOhF9GfTNpCZQzmAtIAYhzleoBnP6nUqtzvnO07eYXWYc4rm2TJdBLs8ncDePOMz2UqlupSm
cGhqSwoqNWmq2Ovs+Ai08V0BqlnSCi435DiuG/FpkWR2NZM6wuqakoVc8bcXKR7mIwH9HULigM4a
0Lg7LcR2oYR9Ouxv8vXuFaR4+1Yq01zZRsRfxE6kjVS1g2XyN1x9FMp95WRcheiFvdlpmZixnpeU
t39xZpf6zoIiJu/sGlrF86Sakr4R9VcUNN2y95HclTtRLPBwJlpg6vShDhku3fBwZO/v3kKx1EWB
z3Q1cnin4jdsN/MEIhVW8e6U/vuorFIP5UJqYHcevQRXiIZ5UHOI/leffHyUDjJ6tksc+yhqNrAJ
krzw/COvNIUwgVdwnZ/YveiezmmvfCiImh7M6Hyk+a8gDCUNU8eoHllxJNAIBuEoQygXcoG5VfvY
m02sz3Eh5uWwoyMa18F3d4qmqtszt/RQtLymPYNGDr/2oqnRiIYaZs8OCNSgyEuv0+jwrx76AZ8m
umdoIc5Ujkidq7BG9yacdDydQxq8uPpu5FFiIGxs3Quk3xTgvjHqEBHM6S9CyGDB1muN06VxxnNY
kY4wNlC7qdvYhbe3e9y9AvrOTXBycyKiwC2tOLZbZKh0yTC+hHJT8Z0Om/fN0w5AcCGMrvfOabZf
q4XFgNqlrqW0W3f/e5y6x+uICIiMa/HLHI23vSlbFGLJS56YWiSVRhTkjZk335kMsyOQ9DvMO9DB
D35GOc4WWdWzqW4zskGiC8uyp7hnO7d43TlWNdsB+zQHoeqmTC/kJnr3vzYyi+oIkniQ6b1NuY0i
gUNb7vRTopx8r9D6Tvw0ukYjsHlIbSpkRxDt5dW61isWQzvYpgz1ZK9gLvbdhCTN+u3QedC7Xys/
EMkp5V2zY8woUroWHvNCXEK2+bY1FYs4JffzBOEgKRgaWj6jzkSKLccw+2rRk+I5dfKaIwh0+XrC
PnRyLdGHi+73a6zmGJtJYqyNZEtY9AsFiniQ5LC934S6zroog82aqvlXbKhdSJDrb8831kHhpNtx
hpCuuSLvmkJQqXFkKdBtmVqXByNOKBFaR8AwqNnQhc6vEQUmVLiHQSp/6/+RahxJGh5W1yF9Utaw
Zqd4knT+iTzEqMS9kM8yDwIRPZbeJVIh92JG2NMUam3el9nYaJ+AoRgHFJYliOoarlq+Hf/A+q5H
nzZfFDZcYhwDBKETs7kd1fZPKF7XQlugQvDzEnFRUFof9be/9Dj0t7i0VctkkoyoJG2oKTSbv6BD
1g3mna+yEE0zfBWQXa8AUD9cRZ/y4Qm2OdyB079ogzbYmaCaPwEq9nDpFj1UjS7wz8Y5BaNhmwSO
KeshT5h4X2/s45tABM+U0xLZ99ssXfLcF9eyUjvpaR8P47duoWXhVSjxt85sCyN49YyMXE+O01sS
FcvXmiPOEOTJNma9ShqA66NmRTbpjGS6kx7QDomCIGJmMNW61XwM2avcjZ5cw2kBrVRW3+gS2UyP
3wtDbvFvFQ5dIvWQyUIBGxV9N7jGPAbO53/s0+MnPI77p+XBn3JwCPo/iXcO90qXX54sUEMbm6fa
j5kSDWiJZTnjYwL1OM17PW7QH5++WwhzqGf1YiXvBnkmpe/8AP4lJJoeOlkOs9r/KqtFXk9I8WeC
id5hOmRh5f1n3fWWQFEVFqYw3SOT38kHhmgs5weGfO3rBslwA5jqxcm19sFyzB48CSMP9JxJzYuc
ebhCJyEMC37o1vNU5bn5FP5ltezOfyb5j/kcg0v59KO5ak/wFa8dvrdHbbgvMpRuOC9ZtF08xk3Q
6nJkyUULa99xCm8oJpuwYhGZElFtytX065AUacKohqEjjqs49L2lTq4Gtdk+CP4ilbT00BKtNnXV
JYCwjww+bbV5MwE6uyLpujZrJ7O2XA4caVhHHqRNclUQ4PLLRhJatx2DqFV8MJII1LtRqh2UvkhX
C6Rj6Zr1Kbjza5zchcxQzuuD1B5iN5YkxaZ+F1NUjv3aLX0Yn7TCa9Q5ZUknTjoDDheZ2uI5n8DR
bWlMiz+scFvRksDlel5TIdnuYkfgwkJZiptEIZ5ft6Wu+vA10h/iZR9ksWsPVdlUkUs8mHgjnQcy
5z843VPiHfXAHlhSMAFsfwYBkFRBwRLLW484XP/1znoPpnKQQ2ouczbqR1aNG1oSDJSUBkiIkG6c
RpuyCGT1szuy9Im3ZBEaj6J5MqfUFfW+t/gDOHJeTX5h8rUIO7zS5XUQ7leBwq0KCkFv1VVKl0+a
PKjMMKT6FKCoACPZIo82MPSj/m4Jsk8MCvZ1McXGj9iAHovIpv3PO7rRklA9FMRfyZNbdoJfwCS6
+fd7j75VUcanwE7QIoQ09LbP5A2EFiQATyQLf/ln550w2hzZHPb6owPvfXstiZrcCKiQlQxIjMB1
JIICMDstmRB8rKHeW7UfOvZuZZWccCuHaZ0pdPXDk9Yij98BDEi3EoRsc2fGerFJdi5VRtAVHCxG
buDAQ9YJILWYiuV8tT62+UNQ1S7s9bqkm6dMTRms6rKpBUdqF/9Be/goXxzwuOSIY77Oh5wcp/b1
8JvyWBog3u8ZZhDm8NDJFkK7eg92uq8qeMT7rnvQ8xNZRnDNCVEykA8zPTwyQ8NkwbH08nBYtaXe
1C4ODcyvMJxyLQwncIPVqIAA23AR4elui2hVrwjXSoFqbtvLAM7j/jNRdlEh8x2Unm7ZIBZy82vL
hQeRZuyKITdb09ecrHg5LfClg00VgWFfzoxTQU3OCC5ZWW6pYw4WHh9GVIltNXhLJSBQBRqPwfHh
OpfDkabVYp0remoTrmQNB++YzdRwhvFqLbTgAbNX1C+Pt0W4XF3+ArkRzB6fxHSltSG+eAn6tkOn
QyxO1L3llxXzYh3xkNcD9ByGwVnsxtGCE7uAw3CyEkTMzzp+kucVR8ablSN0/npvwVmXU/Lammvk
3PDtacTLk8nixESH+AOJxHvHaYUtxMx3doRXOHuE8Ls6GWYVks2ZRqEWJiA3IJtnD2Q0ZygsYy7d
E6MUmEMPvW291uobctxbuMd3AjZUe+DSCvRkB6lbl37Gu+0FDq+2kLysBEjCNxfvk1O5eid+263W
hsiOZO4WUJpBTGrZvuMco9a7fRaHqXEgbjtUky5OOk3iL6AqCgxZw5dJf5NUY0zlDiOoYsCXqyeo
rabIjmPFUkheZnErGhLyHHX0Je+ZxUeVIu0UCosVGiuJy09ypObNUFWmIqeT/fi499Lk1vdjPlGy
0vKDWjFFZxAS7du1LDrydbLUe9PubS5M7WlYUUg1tqRP+ELBU6hcRNkms3GRF2LZYQlGIXJCzuTb
YOJVjclueCoI/L9tQmV8DS/0EEWVyGR7/fedhEbgHl5He2Z7nNX+5TYWDTjU6bYIqCFJFF78vlS6
ubJyCk5Em1cRs8b+FYAacVE2RpJm0I33+gwR1l/O79hP6UC3/SBhscwJm53tCsoqckwG4H9kzux9
vJM/yR0Xtv0Zf4XOM090WdNerDi4GFIsHs/5h+O68VY7Bhiid7tgsCwM/teAh4PrxcewsFElLVgc
uAdom0JK/5Uo6TGfPSMSBwKhSo0jXcpD7ujqQB+hvbLzcqKIR9/5DvpdxabuB1idV+1uNMcZ0M5u
T4vWrHH2XSuYRXuTLiB2cRaByWDT2K508kitMAiYJG4nm65Q0TUKIGZBUMkUtecPUxKWUu17UhNt
jDf0CANvU123SXIOp6GLCNxaeBaRqjok0reXmLbSzsqKXEeohJwU7D/N9OjOW4vq8YViOi+ytUsY
3vA6L3N7cON5YOnpk1pwoYM9i4MnKMWAShr/YKhgwlA4JtHe5JKpeTqvnZq0e/T8GfPxp77b5wt9
Un+IRxfAtt9JhkJ+zc767GyRBKLeFz/sClfBmQx0mLfzWqfwIQau4ocnyW9lBJu7A1evga2XU1OB
GbsmkPDwlH3IbWnkSKXaPr3mP2C3KHx3xhUnvZ4W7jAPwt/UkkUVVmhUmAsbSV5zzIa697py9WCC
9NMZDGIjOuhoyfR5oG8HW2j5f7LLR6siCWeD71fexV1fkCg4YMdHghbbBoNagUcdHRm1vt91tlHa
Ev0ngV6sD+q1Lv0NoubBDqjy/EtfiCVIo8T4kWIDHtWO/YZWKgIwjZq9qraRsIwiFFi1mnA4h2Bo
Xg150prmFc6eYZACes5GFBVuwt34h6y7Ok4sBq0eHgI4yeZ1mB38zKt9eh8rNDUS91HqYDUXwyTc
iYPLhJx30t+V5wJXuDDk3yqj4M6x4hQA57KGlGHdAdDpm6fmcm5FUzAWV43lHE5ZxWBBi3mbjmZz
2K6gxRWrty0tpEROagsSYjy0+V2y80Kf1SqWOT/c3I3EZWzqLMlprzur9aph9/CuokJ7CTo06Kf4
+2MtIiBmiDf4g0mDbefNqLLPqwgQSo0h46BKW7V4nhGkYeZDGy7AcFF9X5d0wx/RZIRfo11ondmr
qj5sUD8WsEIwIj74tDbGTiGtG6PxYc1B5RLdT8AL0QO56EWH/vqiAJ2smCS1Fdra4q/Klitl42YZ
FxRo/SKCdrWFE9S7XlK5K6nbQ3b8+q7WGe0BaX5SVSZKHjhXOc/AheCIst8WPmgZRZp85+SoaTED
beVCTlOQcxS27sVhdiIz+NnTCgAFWH9Aj2xNpq/Uh50ZkGp06gb9SXnKFLyJ93677XNXrw4AZYj5
L0xjBzTzEG9NJiD7LD0itGmT9nUeLTzjRJ193uNIkXD3xhEdDyaUnC4q52fBjCOOtt25kfKy8/PO
uo1TzjqkjYXwoARaU+wmiBfwQHgJ5rloBZXSQltywNbtjEdYBy/cX0t3hyT7k+YF48CFJt3atcuW
U4f5wPc55IIGJwMxISh7wG+PCNCs8Jt15ApTPNGDrxNvs8Cwq01pbc1D7xZmFK1FgS4vjuNwfBdE
PSUVGq9GxyQD4KvBUjT5biiPN+J/8jidil4q8Y2wJWAcHRwMD17Inn6wuiFxU5aiPlCciyfwL9wU
tl7VTV8VFIECn+6LWv0GeOQ+xo75NyxQC9KBnFYOzv9rz431JUvSHd/lulcsZ6POngp/95b2YUIb
daSrKI/23xMZTDIxXZQKCk5u7MDKMbsX18MiymnXdzDuvO82ioRyhfrF8byjHxc6XkEya4pko2yq
rh6BCwLu8zg+aZTurtjsAH9haXwhJCX8vdP1FE2o76tqEx+pj+J3ox25TbdBiQcsIWzZIt1Fb8ke
SJ80VXGYrzIeFBhBmnjRFyRU3Rh7rjXEdnuHAnXOi6NhvQ/98TnpZFeIlJS7h82NQF7cDtLRJAuP
zFoj15+kZ5mVLlznPuDhoxrCQ8VlqefJUjqGHZmoCROwYooQf2Ge/vCCd/UNysKLMd0lfNqCVnJh
ANnNFXPbW9Zg1phKwHI1A6WcwtO8Q6ZkJ6Hx4Kk+as8S2gPepinSyfewm5hhLkNLV/mP907KqisP
YamVfWmtcu8RqQF6xVIqrCp+peQWG9ye648DvWz/DD2g/uK7gBoHURin/pqhX2qpV+DjKU/k+nVu
m3GgGsPe2P5CY+mLKT0qCZLfJ2VzyJ6bUrqbmcO44tdwB12Gc3p1uKyN11/v99H3TIQ3bNH7ydc1
VCQAfBCMu7Doi1Uuawrj3XOYqgezuW02s3pJC0/+3XG5OnRiXMje91hbnn9l0U6Q8Z+TIpIxy1Fq
p4OS4grjnVx67Z0uB0m/SGYwFlvs5hxMnzv3i2g7XZb6AO4jW6J7E5oV+rzseElPx9091R8mHKwT
nux68weSEAfGE1zdQHYQzsVhhybQZ1AhyvHj4EmQdW/KT0sJDIA7Q8AmnrIi6WWiR/KWOpFDtlNc
dAOvyv+C3Xhi6FO5l+nSDzJiq1UcKXENJGyUWH9rNMh57U9ejP6FdmP6h2xpIIUtP9jNcgrbt47X
gr5eJCtLvfgLoIwLgP1xgaqflXmmFCF9HMWQFLACOLz/il+hljQ5Cg6si0C+/C5dtm+CDYOpd65B
ww2ITtxIk/hfFQxgEZ4rrf4tI8tcaUgfaZrsuBhrtw/PbW+CljFEnogSqXar0Rb5PoGuEgm3f6fa
ZcdpohHmRjTvYjGat+jTi2Wja5Pmig5/+FryZWAxmk3U20OKWlvyXcab22zmW8XU2a9TZIxkqgS3
rtFcpO/QNCCBh4KM5pUxbTvqp+Y4FKDrzDSCoWzvO2+476oNAYU7Y/4RB0k7nunTzx2HLc2ybk0s
S0TspjOKekaxIJ05LQVnV8ZCtbPisbacax9T0gBHOZamdL6njIa9WdEI7nPDFvQm0mnca5N8nat/
u5cwt/His+knfI/v5M20Ew66v/fywn6DKTEOad/FKKUTWuhDxcFXW0255aG6fYSTYbJRvrP9qK06
6ssYJ7qTmUnuaN1LnkM4ChdDJ0OrtJZ4bThGcEJqx/cmiKzN4OCkDhFO22xI9X2IEMQudUEKcd+O
zYJhEjXKzOA2rYmno75SuNXG1jyQ62GLrgzjSv7p/+NfCMRBlb6C/ZoCWQHkg4i4/O3d3r622Kxf
UfQmiIEXsFgiOSJ25Rx6YjPbzvykgR9IZJUnnpkiLkl1l5Ml9cSO4UkJ/3XTm/lRrDuTKwk/5P5L
iL1L1xV0UAZslrOxBDoLXCg5aTkMBBgHkZLnCr3Z9MJRrHIFvq/2egpZtkxEq6/3Jbs4aYn6Z3m2
BHWOwhRn74zanPTuoYu3S9Px+6nxJ87Xg8JVl30iNVTskYwnlJ8P635RmZT1al0c7M+btgHEiA0M
4k38NhWdB5t/tL2W3qysqa/t2ufoWjbaizSTdA3ku4E9/Zp8EJSWCmqGWqdC13NXXE0CYMbbxm9m
lyyoV8H6/ENWo+LPocdKBGaCWIgM4afA/aqdSDQliTkzIBufdKfzuOcRKVBD1I2ID6vMLQhsqj/u
qSpuBqYBCUGx9kvWqTDX5fwHv2ixNIxEvu9y79OZ32S84OKOMuGN483FOLOHO9DeA0/ZGgvahiyK
/aqujfIaVO4vxb+vgQ1x1yZlwElSNSB4c1Ov26h00iLTpaLWlBv5SwoTt4j44FhRhc4cRpFlPMQW
sulHlzcGrV853cmjP8LhAWCBQcrnwRe1uGd4x6wE7Qws6933D06DY10okDiuouA1tKIB/indTtko
JmA8hCaB2DPxcoZfB9NuLGqMFmylAjjgTp14ANl5T+qH7nH+7J7zDiWZbDCWYMlop6+Zs2ZO4iWE
oGX2xGFxgiZa0cK4TnujTptXEiVxhzMnR4DeOSsoZzgQzOyCToCYrZIpxqwAKL726zEiRKCUfyQt
mFNbN8CeSHk9W4ghgqYcekYfTEOte3dyXBmk3C2+0xm3+a7cu/c+v/UuqoAQuC7p5qkFRnGI1ZvT
XzuaTZNVYwxeyzMedn4S/racVpJznUSBXohEkyMSolL+FuTMSOTEvat9O1pVdSXTM492LC3lLDwp
W9OJ8XT9ZqHOjlfIjhrps0qc4qhR6btkKNEUJ+amqdnH4LMSUFqkB4q6fB9FF28fQ7wSXP2f1Dq8
b6aT5mCZTbm8DsTj9bWZcQL2UBC13GBb+7DAcAmxzqEELAVsvgxuTb3xqcYciwJsCA18Hcl4ltou
vDF1EgHsSNzrsPJZGTN/gnel6Aoi/w5S/dxM5SoErzvHLJDyxSn/yPOj8C4kGPsBlesS3v4tMO3M
XC+of54RdlhP7o0LaULCIQI83eibxNxl0n3QvWrksJvREKGg7vVUeygBQns5OUePvLaOxRI1rGaB
KNzvzD7G4G/kuoRDIhsfxUSCGTde81WLiZ2CIPPcIRL2JmCKPq5kdLtykwzhTI5rXevj0HwnK5z4
8ss0UK/JY/HP/YSZG5tt/6zb0wC4lhLomrGBMYx971zbvAlTuBxS8BjJDDqQOnOcPt7vW39kRkZ0
shoEii3LOrglKqtw7buJ65ykox7NQ3lrHX3OleVwrPFd5MLRkqB4KjwtHwOTOoNJLbLM0OecD9/w
SxQ3eoAQcQk1bieItOsBhglsr97UyCuWB1b9IOjIjQ0f2coQrPSk54fCA2DHR2OjZHqYNaLfcvZk
OlOtM5loqvc48Jl9QequhvWTvSHhJg0HsfH8PWoda+Dm3ll4GBhzY0jW/eFY6wyIgziPhOHP+7qF
ridRgiMgbyrrGXeUvJq7B6HMI5RAjqEN/obRurzPXKmQLXY/sc4u88ZRKsjZ2odyJzytkaYh89RP
+Q+VG0W9UdDVjLGe5+coKvcK2Dj3OQVdP5FnSSKCnZZdmS7O8sXm9wqqrGi4XlYPiHgB5+l/j4z5
3nC3ipaStyBcXHfL1blSez07xNEZxebE8mqG0YOKEsIGEXIOolxRXiWnbo/wz1nEU5bvVwycfZ1c
DmB/YzGIBxfJu7M51vTz11olvouF1uvOc1J0bJs/Np4DYOofVbSzd0zv5LPgxJRDz7cxF4Lljzj6
QWelJ0cOTHkUR5QVVCymL7BvRUBsPszkMCArJ9MoYY7XAriFnosdWj+jsCgI441gbDYJuTDxZN9b
xrhWNvD9JsrMBmwqyM9AbkoovSFMxW8gZArRsQsGEJksv7AqATV7d/fohEouFe4pKcqw8VHtCbCX
vZEcm/kwY+ve73Hx0kqioARCvly4l2b2nbj6zj80siIuO+PqFlpelDnxkXXBNEK9Gr0JeIy2BaVY
ajbSn/PTQVhDwQf8KbenqToyvunGpRDmxwwg/08vK0JNA8N4grjxCM5ybFh7YejnFwYm/2ZJ7qJx
dDrdakNoMgznI1EBwg9yp3G/yTFqrH3wWSFivk5Ljz8dxyqVOP2XB04spcoeLx+AHzCbyU+9n4qD
FAhfVpPdfSH/ehsce8G0swSxV6lBCCHwnvfa6QiKx/v28wO/A0rWVy+5WmxxwYZjEY6b+HV9gzqv
88wDGjI9vq8zxhh8y50O15SGXObwfGRdbiCfjOlhKN8gKKovCo5uQ73kPM52sfwLxwzJr1vncVo9
KpqRqIvVI/DpuUV/H/f7xMIWHHoL/B1z9guJYnPUT0r3D9XjwNeNHkGnA1MBzP6087p5ZfuFYm1B
eh3eFmm0NogO3k/9qD9IriG5mGxqX8yRpWxIvVd1Nt8gvhgVGtCvtKzLM5T1Z9MnJVxOVneRycbC
BdISWmhfqm4pWmKvMhcLoinCja26woj1gUCAZnyzq2K0yiYtIJMT+J2eMzESyrQYtz4muaH0/KrN
fPwVKWNY2BHjw4bMwwZrr9JTz0uSKceRqYAlzdfF/GEFE/4goZsshTOq56jEgMXoTT2zOffTxLNN
bBLbd07skt+TFC16bMmQeVsMGW2eyMRox3Hp8JK0jgt1PDPq5NRXqO2Lsu0/qU7T6zWjpxLy2q6g
+Wpi5Lbc0ICoPfWy6kHAdqXoehSI1pd4LItsbeijp51fZwQfr3QQZadMRNT3nRFnvhrVJO5labcu
HkjvtfwSgxw5JwtgOWq50s6yCxeVQPPeqkCYKVALXjo3AnC073OeEoqpneFYAbMxgXOrl7RQnv9z
7JSIUc1hAdBzg3afu/iyq9eJ6EcrjzH6EA1HAaoc1ovxUw8gmi7AxmhAcOsicDu5rZuS1k+RYXpR
N8ezNGi+5toJ+FL8a2u0lw64K+5clgYO+EJ3yOaKdikzP5ZJ6pKcgbJMHxz84a/BBYzPRNwMJxTt
kB0F78we3zU3gX8hFpgbZaNDl6OxILqCA65w1sdhO2J3ha/ap+u5yzwLi94Ljwu9VZmRCHUbplTv
ZqnJqTQPNwF5Fg/jy314iEr6Ey+eXwldGfQwBbmagYLs53uA+/5DPJsYXLSuF0eiE2hZRsMumYqG
bOOFS1SxjIQr+bw8bBJw1STkq8sHpV75yEFVv9P4s4bgrYv2NdihV55oSTR/p7SDEHglIo3+9biX
abGCMPqmRJrbMH4fQFCxhe1ItTs6ZQPSKT+qMRXQSEe3ClkofeK1CMDXJQCGddkbsUye8ROY6v0j
phV6Ys5nYe0o0Y1FSXmOMKOUAeVt4CYG3bOr9+xu/zGb6DXPEqv5vxKn3fglLU3u/ki0EXZD6iaA
RZUH/+ODv5D9Wl5sbYgUV9G9nYWouk0JeyVFHkdXpOGF+0C8ZSgb7ddxNvrZrKEvxvh/t/qujd5b
xkKdR+/2f6WalCm5ZY9KIl7tVfHvuSzul3U7NU2Ub7HgWUNqzRg8kNuHjnxdUQgyD40Zyi2bdfD5
Nf5q1lzYliy3HjCwqpCaSmiTWEFvHMz4zmkF9egq6A8XRpcDdAUL/I5fI9cOemhG7yAs2wBi1hrR
Fxdw+o4FMh/UjjDa4jI1wiT7CQEKXj2jWh4M6nQP2TeKQQzjsjpt3HRQpfy95IZcMpBoAXBFVWer
Y1/5gITEEbVStA2/x5bVSvUTnCN7oFC/gZ1rOqfgkul5kxJpYh58ibmIVDhAOqJjwiNZtXDmi6HL
PHoT8G8qdjLEtZA8n9EKwaH5p6EA1TOob69cXp4rhvJsayKVuT+7VRFrkoApEdPkJ+yEQoJLPFG6
+kqz57VHcPCaejE2dDu1qCJD3FldIOVjLw0llUSvywy9xnUfXVbuYCPeyaPMtqvGeXAXuFN+MZCh
LmR8CN9NVOXYogcFNa9nbUcgL1wvk7n8ZM5RvfQHlPPz0SKf2yiwR3nDBsrSeKHaXsO5D2bkzl2a
4iWOv/JS5jLv2ePTBb8WjJEkiTzT9Z/6nyFOCstlvtzNgYAMPzmJOy43FHeQcf2hRZf9XOGF2v1W
uzGHAEVCeHb7PVaVb2UpVmXPPGhZA11sh0neU1sgTPF6Z2LKwkw2gYNYYEemjOXR+eARmaQShUjA
+Sar9jym0SkxMfGUgJxSN8UoXBry5gI5RiF788BPxYvbUKPOxkoFJKujKbrvs5M605xMkQa3X6yv
isecDD0zpXNUSToMPNTg8MdwWCL/ilNV48r2f2DF/DVqvhJUekv3IMH1rkOfYVfDXmLzaGsyhFbM
K9kxGkHJFK5fhRsdplKkV064pBD/2u8CPU2aZi+PfzlPCt6DcBzc5grvGprtDKlSs0bIb6gK9EdK
fXuoXMN3rJ67bnNLPEik7NfD9wDxtRfyRLJqBHsA0mns+QBzwScNgeKialir5xpg9zn4WtLYIJUo
DI8HSVCvZJhxubkxx/dEPKLRUzKjLZDiqwlRFk9J1lWt8zNqE6jU+22BErv4K4QTddgGtbMqWsWm
VVxqmpWwLolbZOVF6juNwdhx08JAir/VqNJtxTmB67mBY/CXSCe9/eep7UahI70nirkT4WotYrw8
UPiNS1tTkJDJ17XPhaif0doL3encTTFwR+WtTl8aK+z/1O/hsve+zXrIHkS6z++Ll1SpmNHaotjo
qKswNwFYsTgh67Dn2PLkqq0+vc5/7kul/vDFQy1z4Ku3GUG0UU2om3VwhYqzaO8kOAjrpyTip2FP
NRFgIolePpx4rR2QQuN7O1Zdt9EA/CtV5bHGY7fJcP336VsmfA7Iyz8+Mw0H3yHc8ZEB4PSj5Bfh
1wwsB1VhvNLy41fXuBJqACjx4FsB0Cmg0PazsLQOHQEuyQt0UUgkSPcGfa2tdIAwonvl3boz9vZS
Ox+cQXv7ylclFZHUgOnt1bBg4mnypyMhS8+zZHyqG+e7H1GXMU38Zpbbi3jEjnUh62s3tYaJwpFv
8505Yw1WaFrCIvabKUowFikXJFH/1Fo/ml1uAuq5Oyxq2RF0sRaV1bVr++yGl8Y+MRJHhzUuWbt3
8kAGAkCCl63vV2Xvu/qWBPpwe9zzJ02H94RE3GmDqxbHKvhUH8s9Uo7FPynC8dtGugJsh8VD1h/1
8PoSAgosjV1JSTEEHjULs/aZUSv/i7gW0hQaE2IX/+cUsOr2vNcyIv5TIz5/eu6IbxWy96C23mX/
fVRdpmFIeFcTIF96+8M/5eqpqY6DnwYjE0+NK/mHm3NeYmZxgx0NVLLJEHEVCjPnDL0l508YpkwQ
mx8AWxKhmJdkMRx2cbVncUnF/p3fyGBXEUqGtFUZd6/crDUzdLfq9EbcWe1VlyzHNu8XlpQVXG6R
2pI2oO1Mw2FCoYRpwtBUKY4rKOmYtKCrmldavlQh/B7w2xWKvqRT5ZS+FuamJHSUf5C15Q/3K4t6
CJqR6g3PblpgXuaIuL3bOZHhEYc8EGO/+30dALgJtf84cpI2DBwwj2Z0v6dsSWJVBo9ERmgEEZj+
I7huOwoWrq6PzhPqrjDqcFGWqzcWtJez7SNJWCAu9MZWiGoNakR34PNUpIfMjA0v9vWi/6n2aEZQ
ls76lZnPGYaEZnlUX+NuiM9QZHFLHSlF032bhUQQ/21LxW1+gp+m/1tQHsyI7jIU2qNjnNstnB/A
H6OA0soGJ2xMbUl4SopZ1UKVsv6Ct16jnoPQFH0oa7dMrPFZYHVmH3oualK2jg9aey1kXTlmZR+z
Dqs/o71O7uu84Y9QVjUMLFciOApsRIefMLFwYru0bDdW7dI7mUMUXOBB5aN+Y2Ryjdz5w5OKxGIu
s0a2VdSm5HgbmZ5rwDMB9KtBFatEdPZ5hQsJjiQBUteu35GQ+9XQ43/qWKyVNs5uGNCXzJaBAogc
t/5R/FXqeWZaNMGmLUUVZC7pGjJfYajzOyxPnaX0AtTKzNZi0D5rwSbVElqrgoW0aQeZU2bZ0vFz
gmq8QYF9+Dge20+jBV8D9hVPJtCQOtzV1i4c7Qsg56T+hORhTUaOotYjF4u9FFuuoF4yrxzRySWZ
RATl/4XEbAPskqvGUfLAJFQhEAJyWXfZYEweCj1uo4G169Ys27FMQuIRx7QSwjQ+vOGsO/XPqIuK
X/UVfMn8qwPJnMHJ5CyxmZgRNZl/m2awSX/PJnVKBLcTgZYQWt7vEw9IwejU1A7XHjWCMZKKXqcv
unlac9jOsMKjPZu+deoy3eXPQXp6EZk2QX0nOdGQG3mTTGnN3u5T8wlOja1g4K0/Sz0dkdPM2k0Y
YvPegKiR12m1j6RLmcbsAsoIG4PDXQYXCzi0ohQhNXy65s6E8fyeoowSo6rxVXT23Ns/+SHZNfvy
AFHBE4BcHlli29QQm59+c4Nce7oOP7dqwgFT7lLGkaOagtHlwYEEFWz6T7+sDmKit8y09i5KcRj9
+w3YPo3ibGjEGon8I+7EhoAv8pLNeL8a9WCvBMabZNLmJsQ3YB92z4PsZy0f2OBnYqUN/yzF+xgD
Abgeoq4Qr4urPdTumqqLzqWybroo9omu4VKvHZw9+lLhPYWIh6eAQtCpvKluDjChm6SRM+exo7nb
R9IgZbakYs9dzExyUhRKo6tUYl3AUH7dwq2cMTGdrdN5IicULCP27JJLL/oyfnPFPi7NgtyOq74N
Xcf+8fK+qHzEZ5cwiNLx7475SzZSB4LvY94pMuU5wUUTlkJMGfSkvm27OUONm67tK+kztF7/ZReN
NRuJcJVUT7xXHzBE4hqDIuZTImT7OX/zrO7z3z/vCASAcWm8GX9fo5H9FJYChUz4V5qoEiffFC/h
bdrBIxBhIKMkoEyT7wWWJzDiSWgARTo5E0GoSMNnLo1XZZnFLVfJl4AuMPAMd4w9CwmSxryB7zy0
cLpwswPqhmZgYcD2orW3lCGyhqwXN6H9c3VuIAueaybUQn/T0dTg8eZqWnqed5PaEjqPMrAyTqrn
WNK/bMUAAIb691Vin2vv7Th8CtMcJ0I5qRnPgenC4CrdR0cVh/8sCOCw78jCSCOnzJPWB/sJGzz9
PIYCBk5RCcGY5kRdKegMXWR7dmM7NWRQ0YWRO+uzogIfgLHqTs6EAD0W/Lz7IxwIr6jToSqG48vp
8VlVZh2AqmTwjGFwxIISER5G5sBxVZJasFXWfpq1wFDv188N0m8mtct/SmQZwoMstgkhD7670PLY
uXPqptZwVUS1g/VXPJJp/ECROlObExrd3TCa/AycDUWGbwahnLQjYkJkPrN+6EB4qXp3Y8hQ2OM6
gNsnvjnfMOnqCdMBf5x41/oeoW8mf0a6bxjvRS7BzHxtkDFqojssas9Tr9GCcmbnSgEJ1bONCux+
oUiqHfkAc67wEEME3f0WlPOReNPzIgS29IwhuUn8ShgRaTjWJ/VD6qEH3qtRHhxsqZ9Z/udVRKU9
O2vAKdSDwWGQlfASIo6g4X8+rkuyzgdpSTIRd7zYiBc7MrumOQPYFIsqR/qKFnxxT+KeUnXK5uKF
LB9fV5yi+170plHw/Dq7PhJdjpPxNTh2vdNk2p9sOEWsujGMz0eq9lh7UJg0iCwfYaYHtq3Gedix
A9KGPbBDFhr0qZdK3YoyECVT7uF+UQ79mDbN2yTno0Dc40/ZA3sV3x5Vz6WS1Th3aNyGcFZcMYBi
KlvXAG+qJDvpPDcg1ntaLwucGB54qeOiW1MevNssOfyFcrgr41WQURp3jZ16yj/aaeSwgpvRpX9I
9w0OuBAAj7qAiojA9rpVszHpDoVx9jYmv2hvpV5uXqOTBhfvg2ZPP0HxqDAVvcqKVPfTD/3nls+G
fNwMFE9ORjcuNBAYKdNrlR6iOo084s97AvnN9DtP1f3oNWVO4/35EIxVCSuHgGoMCdfkbTQHi58N
M/aHf2E0tiSIEIMTYAxmnff1YDvgfdU3SecsmC6rOnyKtalkQHny1e4hSnVpsK94A7KQMu0gyhZE
yDx3zVrFZrS294YgcHgZASaDbyE9vY/b2a4k31vEtCvFKtrrBUDPbK/UUTXKwxbyO3YOYpLBMhrc
BmMJLOQCy6/dVr7HSmYfERUHt/KlV+Uq5POD0jSzoQoKyvrjVKtikwe48uo5wx803l2FVRATGV1I
92BEXFEqgYgWt62WKFIJXCgVmT4l8UW1n2m3nZajBCLobYFcODgUUY0Hc3t4QLsfxscIOxvlu1yh
tr+pT8y/UQmsb45m/ql4v4yvY1OpE4HqV0pEBHF3RKDFuSpWPOMD0IK4l/frEgARaI98Q5DG7uzg
upxqlPIa8ppVUpTadF6J1nK1wrLq8Fca7Lt/WZYgyNrnbgIK04sfk43xfkSGPbYd062jgLcKKkEB
gOrbwdfD3Eu1xAEysUM9Gcld+25jiwN1NvGmyf04GkB4wBSqBQhU8Czv+bnqTODEpioAYMAGUdfg
n009O+5r3c/BCrSwYFtDmBZRA0LpACr+u0p6sW7fOXaX2y2PyK9pGVHBd/M+Sqm6rFdhxS+xbHYw
ekuJkpQyYTOecpKO88kMJi4M1nvh1eVwp4hcpg7d6WCksWDKH+pQc5VGErsowB5WHsnrOjEKDOzo
BFM3Sc630nBHZZCqrBhXdPlKjscsHJ+52GAz2hwxoV1Xg5uZvVHda45l7USfKuYFp66xvMlApB9e
NMGK14AQszha125KWk/jHcK6+unCQcdXNQ2NGj7ymS6ipansyhp1Z/r85rg/m0YGKblUKM7gHdJz
AVEmyiS8kSQpFULTpLK6tOSv6V8eEhef1ziUadN7UJPuDqVpZT4+PHC//NbAQqBbHWTZTIUG+Bvq
viEZPsMTGV50+vE0LuFTta2ocBdzF632VaKKQH5ljCcPXzgpFVSndqXkbScSjIv9jaJPECQ+jFjG
LAkUAhJxnTuUYlLvvqE5t1SY+crtIbpP6Blb+XqoXLfdAVBAWq6+I0MLFMey5SiNH3RBcU/ec3hy
m8h+Kisu8OcsJeT7D3gmdv8MyX4zH9qZExAWICUPecktB6X+nP0c8Mmln+4Wrt+fF07qn87dLWDl
Gxd9D8T/QyrP2WaMyXlK34gDgPRLmUBRUDKd3Zy5Nn/ZMNCQ/zkEFWrZxBvnGJbiF0MY39kgzXkQ
4k+PsJKHaziiXjemj++n7MpFhxtnfZRsiSUp7tG3Aee6iXn8KnvFLpwLqteaERK8IRcbRnT4oYX6
8DwHYkHgqQ81rAzSI8aEWh8F6UuNZU743oNHQ419owywJyf4NvfQpbIuqXsdkf9r/M8HoH00WR/0
Cp3Dk3u9p6+rLpV9Jpttnb2ApjBz7L+GjeAsAegdUqUXGZ5SpAzPSCOjgLogndQeWggSK1n6CXD9
cuC5DKZPdv5WHr63/ES/jKAlymqPQeUMo2/IL9W/I3voGVOUdG+pxldldCVBOZPPCyCHzUN8Yb7T
hZFeqiLwfb3qTPppRJaybslyVO12+rGZEmJtv0C/n/7SoNcTCEm6dl2x7uaxgBCDAQU++5E8hfec
A+C56c0XOyGY466W4c5UZNBXFRaZZCn/3YPpbPrnozeHBpVnpcVSFOHcCjqRAjrsDMNyTXdfIkCh
VVD8ecwkCK7T4xk03GoEwEKFJ9gRcNOZiZny/V2x5OzicjRDcjqZiYzV2xPKc1zzUV98wYUZipJz
0p9wTeAFemSaQIADfWSQn3+b+A+PS6hvwmKtpF1gcypfqNvscFy6+rARpbtzXV9Z/0sOny8r6ljG
p1ZUFEShbPOc773DSL+mtt0UYTAihNswwqyOPKC0E+OMYUZlLlRLfRmEfAKGwPNAHWmD9D2TAPTA
bDzPK+uIFoOA3jOe4Jachz5FAAJMGC6bEm/JmE68Qi3IOAGLAZZ6+T5Up7OJ5drEYSwD+B1VkU+p
0Z4ZWNa/wwhN39uSrxtkJQpsgxZu/pAaMfqaOQKkAkz++/Ur1daAsDVYlQHgJNlytZ7U4MCIwqVh
rKqlMmeYhTHXwbeq2RdxQ1Cb14J+leJJ5ZxGKBvuMEGb0LLnenNxfJAzt73bteJYhzcQgzfthFzr
PDc1ZIvJZonOeC6S4YQL1+qSp9htbAQIkpdSAzwi4tmJ6lVhmdsRzkjEiMVtu1oqf08imKWOhs50
Un4KtvpmCdF6zXwH8qqRux3saFIFKzSEbXzjRM8fxZnBYSdVh3x6QXao6CwtXUcVT+UAv3sjSo9k
HpeKwF1xRONlcZbBHwqWAVOTmFceWUtJpp2IWNgonRHXMTJo6MzDN3uKzQE97o2WVYxV5BZ1YSuR
Tv2fN+aW3DQhu5D7B0GIFXrTBPYANo6G8+3QFUt2UZivLZh/D4jSPViaH75tLK6OfrOE3IsKm4e1
GMI9qnC7btu4GPKcvub/M5STfFlKx5NvfVprOLVOesZpCu0zErB0LlE2Mu1MIL3gu8os+5hmdqUE
DARfnU6zM5vLMwo++ZSnzYfyzmhLV75vC9liduH4ZLy6iPMZFqmkPQcI0n7x5DtOLhlwcLOZtdL8
BiMavbny4atNs91e94vEoNslHHozcsqu4RH1wKupsoKa3LcgFjCOdRmG1IYTIGI5C9Kdy+ChrwC8
GB01H93uSc6KjzGFwiS4mw0nZv9F0RCXC5Zxf/fisjPXdZj+UZAF5H4zuUiao6nIBJ/KPuQOwzFy
AkRCxz4147QcPAfH6VbYff5IHtnzmE1vZ/HNWUaWES8fWm542gBzQYcZVRWZ3qH+T29SgRI1DA3t
fVVazWQgMlyMLzkWD/e0Whjd7xdDVDkYeWKpMsRN8ppMcpKEREqFNRdchVH0yoPMGXP8XnakRNRq
BJe4mgmo/pJxgfANyKBFwSiqojMfn/XXlwFwNIhj1sIyZmhtjADRl/VS6kzo35pzKPHu8khB8ohJ
VQnZeJPM775syCHX1dxzUa0gxlfwWqPSwnCyABJZ8Q3OMUpIKbWdOTEB9IibxVRcvMecs33HXXDa
72XKmb9WRt/yNpo/7whvqmiumNB7PjUnhUJdUT83MVFk2yQLEj/nKjcNM3sXBDiZv0RUumxR+o68
Zu6ZIGaDykGl27rq1ezQUZOpIqqb2KBqSduwkAvwEXJ9lWG+UE1KrNAXBrqkWr7kypzJ5TDKoTHz
yl32mQ7J4MH+VjHPQqyZ7yhh6q4JhfIA13k+bnbhmqq3N1wMgmAJApmoCfy96t12z/wXfbG1GYkf
djP9vp0hjy0AI85gaD+Gxe48YXEuFdq5/uG+Pzc2LuS3suk3TVaT17dP1GbMJUEXgkL90IfjBaNy
FJkhe1/m8SOMVAsl1Xsh6d3aYKYnElhvAeGqpgE++sVmWzrenDMNKfditpsrYOsgEN1yjevHT2yb
XzHs/MPfwgBLe+i0/+SM2flRMBm/YzOhvlmUnDjjBuQGdu3/fJ1ptX3/dJh+hyV49GI1q4fLdX85
tp2u8jyQ+kxtr92VMpzyhG/gKiqlDxkmVINsT9GQi7LrsT2pCIU+nqtolhN04TcRe6D6NHSXliwH
AYQE+lxIfFVAbk6irM4ee0McTfoGHU14HJi8o9i0Hfps/boAipv1gLPckSJQTZ83VX6ETvF2asoT
4UqEp/cSMZlcS8JUzI12WYt1kOUx02NN7+ptjPXpRHZbulsXKisNtXzbuNRqfmXkAqPLHPz5siti
Urbea24mfYzYQSlrDJyjqD4JSAX8+E7OtNhTSQJQZ9cT+8jCK3xFSDve+l9KTe6FUAMg6OEmupy5
InZBmDaYELbfte6uxxQK525c8bloMwCmhPMAIUACYaeIa8tMv7FLrDmRkXyBynNzJ16wkvv1/tPO
R7P9ok5jCbKGJ0vsf3Y6j2d0xCQTuYB9RZqNAjj7W3YiNgeDjal5q2m4tbMUQ+fPnqhXwQTxYz/d
QRcUJTKXtcPZR4wTDkq6StfOUeOIsWwaLkqIuVNwkT1WjnDrG+uxXU5LC0zOb1eR29OJ7D7N0wsF
T67t6wkK+CFmyKO4ncYnQTOOPWYLfQFf/CvbK5nvdlecsDfZ56H+o1nTo0QMRnxYegrAxXpwESQ0
XsAoOXseMrjuL3o0yBeBtkVWm0ZccsaVWUyCaBj6SFNA7cVRPd87dguEcZWrWDmg9bfA4RQMTi/l
0ZQgP2zZvAurKH4LH+t4KTosAMGeH9+Dip7/+Ct08vdUzCgoUiVWPOx5TzZy+4WL5M2tYKLeofRp
IWDAtCQEHzJPFL7Y3ebmacFHvMVzK8KZd7GzN9fkqRkdps5tzlp8oeK5+zYXOrxGRStUgvtw3S/I
DwYNtalIMXjLsVlSpKvKLghAgWYAYKNorGu9x+fltRQx0kqFbGIwx2eOdvOu8qxRznWdk9F6GGE0
xOMD5gT3ybo1c1UVaZAgfHNFbH2OsG37G1oBWA2HEcXi6oFWo6WBJ+7Ff3YP0MDtVy1jSPpftEz9
v1TNmsWGP+i9jnSYmf7jjL56ZsleKJ2iaw9GeNktcNsokENzLT+fv3gWztrQJ/xwEWguRTPFCTIg
XJUYLs6/fa6jIAo5s5jlVTDUx1vkMZR/5420Jm9ak0+ET5HVEprea5jqzqsTYJI8+WLcH5Xb4TwB
0ZNHaFuw+AM2wKRukXvnO+Q38zhtvLMi8S/SpwaP2r6JJn5sBwPoF0i2oPhFJKVP4jChBwPFxPg3
hY7SPbAD0GHPq8IPT3po46AHSzsrqlOl0sihuKKan1CH7/SG9dgnQOnrTbwxrt0PQFcmwbndX4zB
WqepTtecKMr++YZRQtrGEdIrWZUB+kpLc737WBbPEoCDPKN0sVmmhSiwDGlTT5URR6AqA+RleSqa
sPCgNYggog6Ik545EFzFfQYDNBeWfdAmP7ei3uIxdsQQHTvYOG/Mpaqww60wm4Vd62lZEO6ZkPsq
SHmpZAu3DczlczOgHwzaO5jYqCBLdlDcGzRAclKL3s+5p3RFGJ1cdswbA4KrAePvAi/KELuu5w/9
UX9t7y3GJxfjqvCGYg/ABcgR2ZKjF9dtznPfvyZGbnVYNVHEfAwqNF3jtpWGwMfyR7mUpL6i97ho
7oCyrq5/XLV85OYU73003LuveDubiBMUyrRw53lxOmZWm5A8/x08IjBBuj3LOh9mxpEWS/4UQ4we
2baavnW3CYOOQwSLJVgL0MOBePmX6T5BgUU9kzNKmw/2NbBcBKVdi18dDsHiKOVGutLBkO9Hw9uY
m5MbtzjxeCvY/72aPDugwu8XJRDFslvJxBGOIr37BpQyu64g6td9B5Z86Ol9Ik4CP1DJiFwm4sni
gkq3/gHVS19wdeZIykN1gUpyNuaHbPX48zr6cTFEr39e1wDCsYIwEhOoD9q/oAvTCBVrVd/X3iTA
T8XfI1o2GXQSCgsZJn5wRUMT25qP7YhIxva/2GMVPPZdvYZW1dBcTPKv2Y+rb13R5bAxJqtDodfR
3xYO4+qAJ62yD9ZYhXKIhXeaDxwscDCh+PcbMPl7l3sa8uqjW7J3+3CWU9htpw32jn6ItnSdheaL
lalrMgVSXAqdfMqd6q2Gl7B3lv6XWq/+34djx4B4TOypuEG1+e8PS4XWeDOAvMgtKntKL3deUx1k
ZaByKggI+u9QzGmrUF2umaCd+AUUcRR5PA6ZqIEh1p2brWnZLOdgHstd6+gs6YYgQtScCXGobhwf
RrEPtMLJPhBP25eNQJstmTt6nKe5C+ev7CgvPWFIyCTIquchj+v7tcTVp3Eo1bnGW8AY68xlsZoj
UPGrO/l/2sUi3y5ZGRa4DccRGa8GDutyKRKs8GV37zGhKBszJyrftDVMn6y0e6pXGLbx0/9I8RG2
iXeRcBQRbycOySuH8jzbL/tuCKW49WEH4Fy+udTKrOT2GPnv8six4zf12I5OvSrCw7VnI69KB5IN
aY3hRDe9Ey2vZyoawKiUUJ/9UUTGc/XdmheLYVDjqG0B3mI7HrNoReJnLAFbn2ga+zAbsRe+oCF+
YTVV0ggyYLyp3FrXbk1Ty10A/AeWjlekiEl72TVFwi7zGW82z7odGbsvvjYtmg+drL8pKYXqDjtv
hcdibOBQqOMvLwMY16oS319uUjr3IZneDmBiks4tGrNY4m9hlK3wulnWXH8QjG0lPVXcxcioSgRE
w3tIwbJtq5moNMbYf+vuagvb/VgWIFzTQXS63jy0bsm4IyFVc5NusTLpIVGsI2RbNGUsF7CTi1FD
MjfHNdsMsq2lmq3mYY5iCxnU1FhR7b77yCflKFK4eaRHHWGv5+vtwgi5jBEGcyJa4vVHSoObN6R3
wyUcn3OdHvL/ubPsuJQmcQe0tjuuQ7bGZ103ucWldHcJpjviQsFTyAuf7SX7UwrFd8BBRc6kHQxw
S698ewXyKtxxBkYUMiXm6nGrL1Wu+yP4Fr6eaSnujf5gqpKVIdQav5Evcyt6lZoUyvQ7pX6Hp+KT
cpHM+vLlQB5bowAlrPcEP9r+UmbRd8ZqtrNIOJfUUad3CH0/ryVkf/lGpOJKYkuLMbQ5Og+Wersh
4dp6ofIPal0KTy8btTzwVDIIOXyvPCT7azfVWGD5aP69hjwFpupIy2bXuM+k5/vC1vpGI+ubGPA8
rPucnVg/eu7JMDAL9UNkdk0l4+5AIZiFoVViA0/jMF3vdD3Fta+a954l0GbQDcHehNnG/YJBdoAp
niEkZSuSJueF7jFvRDUvzmk3ArSRl9vtpJ1ZulsBoOdJDLYufod7iMRYrUaN180Nru9U3JpapCrA
c8FOHPhlAyT62hKMcJfU2W6CkCCrrSd/1Z8vxTWwMcD30D+xOZyVOepGyhy/2FrXlBKGCzELgyAW
zANoM2njKLa9vOBpbqyQwqorYGa+2IPY8X/XMVm4aP7msJ7JRE8VM1GANlgJHX1CIhRHaufslh+l
qq7krjLu5SGrl+xWhtPsGJjhP/CsWJFUL6WxIGnrzzLodzyk/QE6DsFfLqbxgIbrr8sOUWdIeCek
mwBfxZUeJ0E/u9UJa0Cyw389F2ESadfEjyt5sH6QVgQ2nwMTKvnTkECxv1QMx3f84Yt68DE1K4ad
WeyNNPvk7scpSd97DlhDc5+V71hr1v0RgWyrUmiHJKKkYs/js0sQWiBk5WiEgHPxjIhQreY3VxlZ
HhsxMQVdSbtt/sDsr6vTcW54TvPCqd3LtxLkk+tPrDV5ow9iwNoc8Ea1eTqOW1AS3K4O3esCtj1d
fP7F/uuGJHN6wFmsbTM7s5v8IXZyj5+KVjxtrT8411+Nns/V9dnBw+yg/cl4gIDcp0x6oqpO/bu/
5jZzU6rJEJPe0/aJnGFSzOa68lx1s6HX5PoI2T8Ytqpnni7ipljQH1H4tm21kWr1apMBrob5z6cj
sfAsyE+nyyFkCPBV2QH4Zcnhec7mfffYdSB9BvGtX49rl2wnulNVUjZLi8IoI5kzovPtj+HurryF
b7kkDBOfVypKzYgeNwataJ9l12KZpw+iXDdvg3a9SYy4TM+ayC7vM6hHRDDOE3tWYZ6OywO7xJXA
JG4s+nMYNhILkCqcUx2pATzoycT+ZF5hFee3oQ0L/u3c99nEwJcmIOejGZI4DdYgy/WVGPprLp7N
RXEoa1tZXxWrqDHFoxtuaKIpcb7CKnixqeG7hX6mUHrnH9XWB3J+6dUMLWGv9zacuO9NeYrXY84b
Dr4DvxvERlKRzr3nDUDAGAZCK43fr5WzKM2FFBeaEEvaP+A2CFnqqudqNV0Lt4oD4mhhW+NJo/2H
FvT63MwS0mVqT0zwpMzx9DOep7hJSU17c4pFe+XmHcpi+p47dmSmEQLGwkUbZ90VDOxW27Kv6SdR
Utovd95amyiWM4xQL69VSDfwQOJ1RZRi35/vmiXhvFsABJFzHTG0w1YVoCUNCjo8nqIOSS136DW2
Fdt2TtPeGh4s3LDJ5xwmSU/D55yziV77UkrMi0yVO+2utBA1hWC28C5SNk+DFQNfNqRJgyBl1r95
GS8PjnrUjxw4t44qf/X6Clq8+dKQgmfk+d+M5eVDQxvfnmRmcdL4kYir67vFznSHValc3bgqB43D
jnpE1OSKItSzQXR3GEwdDKlr4vIu6ARnhj7c0WM7fxTkhmTHXPitWPE9XolqAoTrF8Y1/9D46fdw
d5Kc+Sch6gTON8DcwB5cwaNGMJcbh/ZoEGKnO5r6/X1/rzKaB3ZeQwp3xckAeakuDCOmMMMVMCtM
/DS8b6WTRmO5J6x8VsseS1n0IjIArnZT1Zb9jGoAMKTxjzIlqsXSLci4E75t+Mu6Yb98/n5HetQc
+TKHZsh1Kabv+L1XSpPj/qoo2w4dTmktwgQ8LbFIEou2ImJLc+fGGltFD7sR/ysPBtFcTYn1dDIz
0KNj2GrVFiit0osMuT1oLJAW19HpkxT2uu27tdn6h1jFa/BFV3/5T6LbCHK6Yq0m1/WfOoJ6YQa0
BXBUXRAdHw6XpmA3nEp6fWL+A6zZr6XkR0NFQcvHb7t9Tj1mY3qSOIS0zE2gco3/SM+HEMYikVHS
a2FlnoPrRviiT6Ezt65xqg7V+dQGVQj/AZ3+dSlRCaeZohDp1eTr+Z2fdEEBlvDvQnlJGhg1wcFP
osT0eTP4Ki/mYzd3ZdWS1lrXJ+W6/OdQgEmDAvDoOGOCTC6rVsIJbX9JD+ucp15sy7SxlnkqdLrY
d0IPcC+3m01i94VcnRilh8pBSg8rQ1Dvg1ihKUQ1m21PcoabkN8pEiMWMpufRGuVzBe+lzpYwKoy
BMPU5A3eJTxgAZ19EQXIbnJP+Jpcc8nEoS6nu0xvjozqW4nkS2O5pmbL4v2mBhjTZi4IkP7SrGZx
gt3lFf7eqfqbRjjQFvisuEir2yClj6hBTgTFJ4iFtd60KrUpr3N6T4ZqdDGd1rqMs+oXMDAdPvz9
3QNWwnlqOK/wmR15dj2fN+Pmb/N+WYq3PPrZEZpudxPrJHRML62W9D1eoKi4a26TEyyJvqIYleji
j37CpZ/HSkYxa1/Ts3T9iR2MEEOgQnODqztYxBnzswhNjmzOIQzwfQoau6R5bob6LyN2lMiE8mRI
SoqnBNSN7D0/nyXKwlVnraHWZSlMYub7/iTvVFvQpSstWRxztp1Sg/WxdRWHxxThI7PTiCFYe3zP
XpiQLw96SQyidTjCYv5+LOnRQcEn0e7X//fz598Ht4G9DwmIHg83LwWzcTbPDMTp8wqhjen7NeUg
mU2DOD6Nh7KrDKDjZ/0LHTQy3God2zlcZWM+ELLT2pJZqDUwWlBzKapLWcwB7J/xQmY8wWs+tzYJ
f+G6S8NPNNrjZz/CRhYE+SV7hw9BKANrwQOdzdJFJbd5YFUGhc6xPVwcHxGW13o5P1/pwM0sbz4Z
UZ9z+DK9ddGuuN/QjGpbU7D2aVtsOH1ZAZOAoEc4enFkA00ozt4nA0DGmVeQspWP0uofOQTG4RRe
MHWAkY6j3o46yjhr/GYjsdTL4uRJiHbFrMErHdagj3nnBNqSi8MYayowkkWoHw6q+P0ReXu665Nh
sdm5TZcMqeWM6N0MaJpvZb3/biOoofp682cuITV0U2OVJ1oDT9fLFrgJDBWY6kXKHH6eT8KfK2ol
VWVC85u88MUbnMbFKoNv0uonTbUFWbJVrP4chracRVHnjSnmkUHS8W2fVPxBxgEGcgj7CjfwX3T8
AcY4L+CZQ06R5tpyqXRoiz11TpDXpkZ7jWryz0VYIdJ5A8aEk3Pb9PjF8KDU5i9VuqiP6SeD7FBf
fAQF8JEDfTdn6nB7MHbRy16oQ3xeoQ8MRY7Aebo8fmIhmvoFUX/uhBa9yiCrzqWlPR8MajrExpG2
SLrnmnbs0YJ7xrA3mywRRsbZDxzZ9HVZMvp36X2afpvf6aTNvY0pQJIWiX1rEsMGvNsLhDWkwrft
TacQJb2YEUTdXfHiOKKY5WPK+a7xpBXTmthDhQm6+DLAnkinv0V2XwmVFOw2A2tBWoIetdw8x1Ok
2ecLy0xo9hKt2793liRoJET64Ny9ELzWpihm2xf6ZT84NHekK8p7mL4nPAth6OEE1HVCnsPmxtUN
4lqUyofVLM8K6u+ZaxiD2MOxE3Eeye7Wsm/AWe3pm9oZkriIi4ABv/imNKhwOtFo/LDkCFDtWWZt
ufeQIIJPf2eln++Ox1JQePgtJdDOte60t6Uq4/BFWrDOkFnI26mjcWAIGloRDtGBhS4JuAEozRdl
VhPPkMnnuXAFwbvCxNf/Zq/2+K+6XqIW3SXKgZg4/UhW1nubT4n6Aqp5V9mxK2pLOHIXbg6uBoOI
Vo5ndGo0I623/53UtqHRatWpZzvDG2q3l0eRtW94FJlmd8RINZOij8mJ0iVHUKwdvzHl+IN1doCa
y0rzEegYFmf+3/aL/QL/O4WVz04QIVFYeZZ9VXAD+AIK9jepVDHrLEQr3miRnBH5fceu67cuVqu3
rvkcd4vkzoXb5Ix5+xqGRqftagHQU2OXx00c6HxUDCLwU3dvpIsyrRDL8pdlOgw/8CM2zGumojdt
5pZFDPn4Svr9a3Q7s5V2i16+8rjO86LxB0GXDu+iwZ3i47Ao6N1b2zve2nDQ3MhrzrhpLsemdzR8
/XrTyWSCdQEIE9AJeahaopAlrsEjnjMJ+dUbhjIdZ9sn7ijVj/Gchuvg45TUn4rRUcLAcNrjhtgD
ER3t6QE8VuGU9pSgTuSebCgAB4hUKSHEEudIzTaMQ1oUABty8A9FUlPOx6/WSnMBpHFOP850XBbO
QQMxgf1w8CzgTYlom1eCC0Uh6LdInH6/Y9QTcjXKicVLBAiAeldNixb8lAs4h6U2Gv5RgyzlGBlE
ihtEBqNslH2JZ/dSiaDkGC3EBFyvKzPGy6MyJH/WHHZd+VAG7c6uhNUc/Llt6yhLFFy41ed2utD1
UU7s3Y9gQwGnoyRnRQeaKhiJ/Gn9mgjQxooVl66sDxmymx7hCCwvfQej9c2dkqDUFvUIZIm7J0EP
T2ABxS4pR9lDkALfa8w7yUHtSCKCxJWQuYZToj62ynHl/0eCVG316254NzrOqxi5dbqidM9HgEze
hL8Igi2GwzWh3XAxpmMg1VSEcNRc2QSfmYAX0OmggQ0IayWbvFfvTiqoUokh1xjpikKiTmEqClul
2uTebGQeZbECAvQmE/0Sz2ytVJ8nA6OeCh7kXOBk/EVGsKtn+ZXlqXvRIlIsdw951eL/uGYEOucV
HUSkjIzTAl9BAMTWE6U0lMEGBnxpSFLUATNLpY22v0fb57FJe9TjtHHtSrT7czKODCTwU3fUMs3U
IYXF+tQWN29GakilODDkmMSPWG5tQvz3bcIsxegzF5EwCj7LsRMUtdL8mPzdsBXnzs/SiJSQLufs
+yLx+vzf8ATCDtm+dfCKGSIHuUjMvKmB/F5VAnqJPTonUT2B1CmMc2i8TRBA39SbFnocJr0l8C0h
X94CzkZNBkxflXafx53dLiVeC/zie6fl+eO798bFtwWUphAST1a75/fTNXKzSMcwDMLB/h0O+5yo
Sv+Q7rloX8svx5F9YGrvANegytDsBtSsgLiiplnBTfzG8RzHDdrVlwKY0adjBc7kxzoNu8kc+4sP
qneDuwL3wmxpYTpxujMZoVeYyZ1wu0bYKyu0Pmi4NsAcsF1JTinFsJpmo7r+COy0G+gw+D+b9sPA
SB4GGDR/9kSaJX+1UrzJiLuXoM4er8MH+UuJFrAfhNQH2qoyUduZ4G/xkFw9SYr0HrKz1kicq95u
Bs1VJF0789mbHfIOmne2fssrvm6g6b4pF1jZzB5dSrWisrx82xziKocwsKvCvO3qK+mDGX61V38Z
WahkRWkhC6AN49pu/gg9v3qkLQpObaqyuBhAQW9CklypFZMyVUsJlOEr+aBoh6sl+a6Ze5KFRsXB
aHAY6jB9hoxEtzsrdWKdNCYig0Fdg367R09djSkQD2WU3BDvm2P0ZqqLzy+41+ZViJ88P52zkxJf
1ZtxDN0rEep3bzUd6IalMLfWAJ0dVM1oVJOwHa3SYiTLsT7bmMZDlLKQn8TpfyHpkWeeqVm3/3Yl
SfUS3NM4d6BrQO0/RdBSKXGXeVWkp6Q8d4eHeSzxxP+eMbo9F0axBCWghnuU07kNWehkaXjme7XN
zOgq0ITk4lnNEz+VqQzz8cW1ByzC75BVPa9yhxFc3cgLXvMcWzalzUbhhz8gkBsz8GZVLTwkcivS
UUXACqlN4VphIG0uIEHpAfISKP+ieDYzCmzhT8L3QJqsPu5w9q9rC7KwDTXqhvm8SEe8nZ1fMWxX
504RyjeUk9Aq4vpecCErTgWDS1RZQeI1GTs32mBRExibjZet5/IQclrOlaHQuLTzoaeRyOCWjP8c
zIPsJKxebNhkK2KqQb5ZZywGY4DV+CyR0LcPo2okia3CwO2Kn5vsHay/Ym1Y6I42nMjF2zRlBhKp
s7dFjwsIuV/oZ4OccJ4AeWbSDvFfleX4HotDbn+oeCvEjaY4GEsByujQ6vO1IdS77s+WHIUyw3uM
O61snyYrUhYBtjgaP25ONZ0Sx6rWVhS2Z3Kqm/WtqyljTc+8APzRiyg5qLsrLfhuWgWit9jiJwm7
KPyV+kzjsv8eHtapUzBKN5iNMBDzJVHybI5uj/zogZ/qbkmdygjVc+sLCcc+lb0I5oK4ZL/0NMPz
w4Sgx+NR/apvK1kw2OZ5vLR67qGzacoGyt9yipWu/zU2nE2DbJiob2a0sVbJNKzl5n08llEL/I/L
Vb94w1Ek9vyKqPDvYWy6mRbwFA/ruAwdoVYQGVJDv8jl/vjyUCKNGgzsD6yKdH4ad88AQdFPEcLp
qE/k31ytpcKQ4tWgaYWd1nLI4kCbKv8Zt1oUWBxSNgB5lrPUvdC1etOFzxfNXKpvnYfalqLI4Jht
n46rwN1JIeFtd4NsGR5HF/0bXrZTMizvlihS/aGlN0f0LPNHiIMIlj9e/4iRF12x+TdNeUj8c7vN
1l6ZXzu+yc7lKTz/EmwRSnk1WCvkKjG/o1IzsubofGRekFM3iYcbfBA4q/R5E8oc+VKaliCLZc3X
nwMfOEzYti8cuW07Px/AvVJEh/LkeK2RGYXbC1jOstI3Xm0Wz08QXTIhNSVSVDXCYlZ+ZrW4prWW
zlRJ0dohVrOG/H8QTISJzhxaP1Rfx2NkfCUWK9Is2mAHBuWAPi1J8t06UBLOTAOooAdePSwgwWTw
wpdIU6yv/VSpG3vsblQpQCvfkJJBGixBpezb7qihdwobUwBhgt/SBRYJ2W32SlP5TE1jnMxWb2IT
pnuKn4yZtoh8MON+9E70E4JAgyqPqjFg+Q69YGoROlzEwkrTlI9PEAvE1U894DfW5VhBqTu9F3Jo
v1LecdP3s0LZtjDztrmPXYkEneKkwY+4/N8dQhtrSvIW4gUjmx87WFwKUEL7vPxAlmnx8lGvEZUw
dVkS/HiX+rBAoN0IOm2fyjThyPfxkxGKpfjwzuRzpvDJVCer8ytNYPRevvQ3HI988v86GyK/BuXE
j5zkKVk+pVEn61lDAporqTI7d0o/ngKkUlxpCmK3tvpyiq46QC4qlaZStideL7s+k/44Qj8lba25
LKxvUhCRBtM3y7Vn/QNp8/ag8T1PFfD/gv6Y+eOW4fcnmuKzvq3PrRnMeDewKTvWOSMAosnjOGyh
h42t86Pm6UWTeXheLGku+1HBBNBf37cCRKTqyJ2GU2LTzTGnmPObIvyxBBXlQjZS64sc0Znj6hCc
jFh4J3q2Y3UYjvkHd5RmhONP2nyReAsW6bketbhFOnm4SDl/lF4cRRkG6HyLBetQ3Xo/oY29hxaV
D2XkTyIAmV4B/CfC4FVPY9OLgQ2z7RTXsxn/NjoNzzJwkdb5hTmb8isGRuDk7Iv5qp/g7mxlZWny
StZKT/nkdoi8+gxXj+bfMfCSEXCXaXqQ5RVJRRbEiy7m2kW1yfmGdCxHUeVHlxg2x/Mcr7IlenxE
dhdtn5/kn+B5raKkVP3SDd+1mxdjMSFVPBsKBaVhEco/nSCYomAQXyz1ZVOfAOHr2DbNnQvvughv
fqzqXxid+giw0yDovJPRI8Wp3f+jE3M7A31YwnF96bCICtMGqhY1+zHn1R+QcWDSGj8ErQpRs7eq
mt8QqPzEfe1uMXeqFOfSGiNUu/rJnDclWtWIaD47D8e6R6huc2DPVnkLgPAW78kZUZAr0N29C/ja
B8TtI6WzfECRS9BDUXEJZdnS7c4hHcf2HObrzYE7vmHlaTXfyrQVPBBZchfunD4OFkrepJqj6xpj
MJTGSQruQUIEvB3YUTFi5cLojxQRuI8+QnqpD5cFdkD/ToEe0KZ2U6I+30j5foiDppMJv+M5aT1+
JxDMtgrK8yWxUw2KXvmPghesm1A+K/sJVbWLEp8zIZaZHSxinV8znz6aNTKZBdWeS39nCuBbyKj0
hm1Ahd5sFrC4uQeY5b1IpKqoeEkAaLVGIcFCc3k1EIGHTOQndM+mWCgnQCFrd0U9jfPmVDXKUUUD
hCnSy0Wi11wQGqMr1oumnz1oKakomXx8GRSl5WBrUXTQOKhp615KUkvtIWBUTzUm4UOTekBKwyaQ
OzS9dcvjTJPzTgXm3MGVvCKmDvzey5BLyMxHiQsJXvZ1r6xf0wGfPnGo4WwlQdYwHFkWEHmSHooT
9NcjrJY2FjEo94K/Mkj+w77kwMkHAw3C8t7gmNOGoy/vPQN8FiVvdnRXIP8pcWL/cbtY2EyUbz3B
2t9iV85CryY2XSjfKdJpj7e1umn/BPCLxP6nrvjzUNx2HquvLlpxzqeZn05q95kOdkASj7cAqtnn
Q5X/uqrj+GJbq9Bp/2VUX4Wgyc2ohrOzD0QMBZEy0+sKd5p00mDibsx7VLo1yO1pe1SpV2E2ueZf
fyNaorqb0Oxwdg93+ocrWKsAt504qAdRreSYy8YQgvdzrzMWmg7IQ7zJSRm1L/kMfTPGlADhtJ5Y
XZhQcVZvvr3xrkLtlp5eU9YcbDSHGMWEpuIokzyaVL+Pi14XJjBj2aIzdYC05GP6+1ILhF/R9XE0
Lh1yZl5asHJnsDFKBjCxYRDaBuiWt83vXh1jmz2c+4CGR5l8bBYWBXSFCttBuMSjSgHu6J+vWhX8
GLHT4A8AtUSGRTLl1ihVR9yQ0LWbVkmoGnwnrKglPzdY1uZmrIPYwQkc9CL3waw6PlHXB2AFisWw
IBM5JYj+vpPPvNeM99wkXN3rh/UmFescDcUFB5kDmLd84FubEn4FBWMe0W/nOtJUfiAGSXqrmyYz
kScFhwtEaWqot44YgFtAJwwKDiRJg7VOXMV4LBQlltjOD4KpSbkN5SQrPiry+P3wD7ZK/xgaZI5B
pj++TILWNY221O0te/J0yz5n6cc8SLTAfbhGsG+IsRuvtGIqTl5J2V0t5X9KHGdc4v+N0r/WoIdO
J9ZWehweZ1TOYbysUndZlNvsPVGaNSQ3zuDxq9KZVMjj3oQRP/4OMGNoHjrRhe8UwUMTFUtMIosI
uPWcUJx4ychX7SOewQpH5iUVENJWp+ZDLwbib4Kmp6UDtvvxWDrjKtIN3sxLDXbKYQrHyRKcy6Et
TEtyLXD8zS73u6TCnJE+rBERhiwUGojsW5H+BFT6IXzb+oJzCFjLoHD7P64+IUfRUHo0rGJfZo2e
4malxxWGIRpBLBLNxa/rm0bE4VUuEslKX/nCuZVkwDTjr5YF8wwZyIJQ7rlMJdzTKiXyzTgUAevd
fF/mhM0qEq1p9zIh+0Qk49aTy07s0fynHIzEr2jbmd6TuLDlqy+KlvpjvtNKFFnjsoG/P/AZJKlZ
kAwnwyVIVwZuz+Xqz4+FTs5AxAuRTCls9rCuBBb23bX6HkfY8GzEJAKZ9dw+THEjfPG1kqafTC94
5T8J+nq4YiC0+GChCjV8HeR+6mCVnqTQSZ/qz8VJMGow5nPukerTSP+uAlfdwUm2Mr/+BVfARpMS
Qlfm0JIh6clborQJm5/cjit4Zyz1pt+TL+Zu7HtQq4HzPqx6URL5HBcw+rHOJ1Qo0Pp5O0Gx2Jg1
3Kit/ddCA2bLuam0uBQN5tLc95gwUaobkH/L/lf6STx2u244vLSK2IHesKTgbfZu0bds2xHPckJL
TpOWqxLK4brE7z0l51ShOtrqg415BkwzeV9C01fpHPh+1kjNbm8TzodfQnhPsttf5/8pJRAjtK7q
1MO4JfD1v3H64XUiBLy7BYhUCuuPYbGItQx3bTtngoUemQVcuMy9ip9sS7di6oth2uKcC+v5Ny3T
6kMah2L5fwu1xobsHSpnffiep3TDlmtU6FzO/cEzicMupd/dvsaFm5t0T9L92tR+E6Dj/sgmHagG
HNBHYGkeD2BXR6/by9fGISH07F93O3aVM6hG+gwesL+2Wm2wawINRXU/J5w4gMky0XFSPvSrWi8B
Ib2UU4KAp85eea5fk4Ei+5P3aYjT2qnH7hkpkHypT1kS78GeAEn+NvE2caRXVlHbVtewwZAoi7GX
ZDFlf3ckd91IzpKxBWQ0roQNd6qwtqC/0bcIGrvjV0kUS0NBcIHfXkNg8/zdIL7gJ6IrpsS7EvZL
keJTmCSAx35iX+KhCgO2syLhlo6ccgQBfYm35+SugKdxSKydJBtwu7fEYZ4os25l0oZBimz1qywK
rkpKDsAnCxk3D3ZMnYZ7IR82RynXIo9Nin3aKT2rAhY4+rah3iEs52s62UM7j04Fv8mHzaiYAxuh
IWLo+PkY4zzV8YopVfWTocrv81OnkOfGRSDFR2PGfLaetbBPkVEKBzJiAEcr/5rb1G0x0brir8ki
LxNml8ZZASufgvDsuiehLk1r8hWR1PN20aJNwAI8mbybMxGry+uwNBOQ3FBI2hW6SMVsqXf994+r
iyffS73sHEtGtLrEVNKKw2cxHjoOqFYwiffUzS95qF6V7K38anvnucllgz6tedodTG90qRhr5VgL
W5Tk1kGrc8tJvw87l/vOfgL8sR0b9DzLU6F6myPMUA9FhRFaFQUFVTPyfPE/tvgrV+cKn58j7YU/
DIuiZRvqslPs2Ma73T88+GFuvCGFdriRU12FsEp+AIU4/OQDa6Sp1kkI9yLN+m9EA4MJVl89ZXcu
kaqEANqik5lBn51GYW6njNCwVQc1nd+nqEezjnUq0q4C6EEaBU0LIhJdfLh9nhQ00dGMbymquSwJ
H0D9/JnFxvQmtKGrCtKIT+MvaYTiepNxCeVVse2QkM6NFHF8wyk7ppZck1knu+1rmzU0zI6+sXxE
Ngc6mOy2oqeVT52DoGCcA2a4zguJoKFnzzgXr00m3E9n9RCIRY4xkmXyd1lr8UGKXkLkkRm8JQG8
b+gReYR6U5ts5ZOG0O2zQp51xuSlMd1GzrTNY8RxiIMHECuWjKt2RWK7ZkE0OvxoeBW7UuorROwZ
20/eaCM/bgYyFdMDlTkN/VUf6xeL28OAklCdLfVlftphgZDJeX/N5hWcFA0uzBixvlWCrrrLl612
TB1Kr/X/q/7Zo13wZy6fI62DD/nTo/B++2HgmWPIdqHRxomrOS2nD4LC+bDdGDZma7NmXs6gkLsd
eo20kXD0J+/u8HLhUaVsd3fazp+ESfqFc62+SuJjoNnki5+WJlH9SEb48oHoV02mqQ3GVTygrE+v
FMC8JNoA24cA5H+PnTQgnQKq5nQC0QlVz4hUf9L6sghSUiC92buuJV7J4hZ52uw849EAoYrEJOf9
DAuGk7/12J1TdOoJAtnMMv8mlBdTqaqmLns5g8oWkTZNm9UyhfydgAi8wwCZbNv4n/QwP8DBJkp5
DPFh8W96OAEu22t4L6nsg7siCJQViD7rIWtn6csfe09GlBKty3mDMC9fAWx9B8KYVsEYUW0ueA6V
hijiL+ce36agzDEHNGpwT1PGeGuhj1uN8Ds6uvph/fZmWV1zcBhtXKzoiJYu5nVUSprBzD3x48lO
GHiZksQg0PA+NPJ5XBeDJDf0SSViORMM2k+4GNUVjCR8VWmXOPQuviJctQyaUXW0zO3URt1L9sDM
cUP+5S4S5h3xUcWbDTYqxHWsyrGBNyORUdpeUV0IlvV6RcAerLXyLv4oEUvxzwW3bA1k4AooBpAw
vKXaVyfEzLo3MLmVmCkKDgk7AyrSPv74Tm8M7fTLTUZVtlbCJiPKURJrqo/1fg4vQdSqDxYSjD6j
FxDNEg1PbHwg5rrtrK+5B8Vty8TP4ZX5SFyJ4YBgyyPTZS3u/PXLKWAfQonwrYZQ/g+kmoOymHTD
/aI2xAmk2pc26jvWPJ6+hYa028ttYLyKdIlsD5ulGrPEp7DUQOeLm4aC5uee/WqkKj1cOhmupCsS
b6+gQ/YnfD7+dNWehQi2F9U2dmaEOP0wtOnolU1xix3B3ID7fYKwtk/1+GsV3X4wA0AgBZmr8Zjp
+tprdfTT0HLdNY5lAmkPKtmqPph84lkdlroHI3+1TeVXPR73NCUZwFZuAl2Kzl+HrY8BXRbUgtj5
CUPSgkXhbzzpK3NC8fDtjR8coBhP0P00+rLdkjeJo7/X1v+drbGLTIVqOaH1KMRjLFdQZz5mTiAD
4nvYkscVcsJ2yG+MvTQkl+HWi8tc4PK3caXYurlZdceMAIWDolXXEZM4mqCHumbeVFDv38xSzOcG
Oi6gRQ47ZWN48CmJeg6r8ygGSkPD6ic1OpmYwMW+44haAeK5i751d2EVWz1p1PbfJadcb7O0Yn8K
1FVh6fleg8rLHQ7MAW9j2WOgGZCjQetIAPv2wBPLhy7DWgKLdjWPkfutvlTkeg9tYFc8tYM2+LAj
3UBwA7nkMVQyltLvv8HLum98cKcLc5EjvF1ktFYTlH4T9+0OERplINTg49dzb7B03EaZlzEL6BMu
15k1xrqI6wyBAs4WpfjX9GUmCerYlvljHYtriwaetVqagm2jzd1Z9OigRCxuwz7qD9ftfAnt7Kis
umNkwwlJqLq5BTGfapZa46WLKjJoPvJFR66/rxZb3/djkVwRxABKAWuCnRr6EbCdN1qdmFPGXKXb
pPyroYivr6teU34oCqvSCZLNJyuId09UQ+QRDe5Guv/aS22H89hO1PHfVxbCxY2OQPdUxB6Tlob8
GeBIz7SmJGDQ13nE3bFTPp1lZR5QtzUYdxpdwiUp921mecV9Am3XCh7tqIV4Hrw1q4SfKaWJ5y8T
KrxcdIaVhL+iriP4QjoLjBX5hmpswEq2hxVz7JdNZ3W+gr1teo8nkayiPYbUtZ7W90xF/uH8U7ez
6alztfq7/mxBaXLKzQST2V1TmNifEC4iotsRJlr0Lwty4ihzx9H+02QdkOYLBWF1Ayr/ctrUkX68
DGyNcrMtqmjrj16QSDCrk6O2ORmsWQ5zJcvTRt6qt42eNDCHfBlfinPP8H62ESJltqaKv0Tjl/F5
+//4TcTqcodHnV7G5vNEI+IrMQR95qoaFX2PFzEgDzsrMuG0E2zQ1E0wCCi66iPF+Ksh6/skaQ8C
CYN2wDO5L3JEsqReCx5Phg9eCbeQqNAfzJhuRpvKx+wx59IV83LjD+50ggNApQK9fDsEv+NGe9ZG
Cd2IJnMexgrYHhwruOwYA6P4owSax2N6pMJ0W/LsSmN2Tbbdo9aFIBmu9XwyZqTqvzG9WRw0VpUT
PlL0i7zOMW9gbj/QPtbg5idiIyK194mZQ4tqhpMh2ZmFW8YTFRv1PoDHhdsOoWN3N8wmQt5BAKkd
yd54f0cQZCQbuGkigj2WBgEmbQ4bMxwTO9ZiVQP3u6FN/l7HCUvPGjAUY0VvIzfYUBvu36Wc4NtT
6tK8nXN2/H3KNNKOGfWUaPUJRI0vfCxypyFXBNoMQFb/2kBL2pdtrvBb4zbzZP+No74NRt6egEbQ
B8dubuV7IPV1P44S4B0kCHhLoiUMuDXs9q1lJasGPLQZBdVgQcV1ZaoPsAKmLt4VXryA0EOB6Iuu
QVarTWN4k2H8yRkcX02SvcQ9q6teLwCKs0cAfQpZRSy35plSZKGjocHrwx/Gpd6dKo+ntYDjSlCD
wQh43gvdxo4GljYr04cLJSrRyhovdVcJlqOxyZBeO3xkFP7YxJ8R4v7Ziu/Li/bfgWXCfcWW+zQy
DD3sROWKAuaqSxixRcmIK2U8irSk14krCwuLZl8xb65/0SLSDarjYoPKnhSOUlngAEdivAa1fh5+
EccJrCTHC3nRAx1+nV14017TX+GfThbeocSQqq1RWICd3RXG3agUDEBbIIRae1xc9G6xIGGg53EM
qUmR4qqIo0D2M/HTvNl9QoagEGW2JEfpu+xEWw7w4nr1fmXUPMlDHjgtBNYE7PbSidQnaCNi0bB4
7AT67PX2qLhOxnBl3PE34X4KP6c3C87RIkmRctXpUvcIYGR0vQc4lAQAK2IbF+AXDUJfO+2aokk4
qOxKDaer3h1C9K3IeqWYPiX1bbIUwXH6PqCpYCF+BUlgXpc/nVTVAF5c6a4t2O9LOr4czWooL1F4
AdHAf+GL7tkPJzEsXF+l4JXYp0zSUqJ7Q+MhQXVx/rGPhvV8vJVL4HgtNLgEHq0LmFPIR1k5WVpN
XdZjVm3ipPDH56u6JdeLjIOiFgwSjVSaeASrVJYOx6/bfO0ApiK0HQpVU7sfx2swAZPCY8mLZXSi
uY2ZxxBCZUq03eZZ9gOJbrMnHrHsjWxJt6O9NDATASxKgU/bHctjtwGf2ayV0vzU+k22xwO/MScC
EoYuLSzmtiM1JZw/yc11KIIn7rMRd0b9zHJWVbMlrEk/F/YLhD4+Vybtjpsv2TpCtK8recydJroK
CnM66UPzslxhidQgDnveA8GVxaoyisobOO+GaNiQ17u4dVvgSY3cXctonygKiUvrXrl+Ubc++xQW
nKR2Bni6BO9LZjkm8USf2lbCZUTwEIXWkwod++cP8uTsVneEAEx2mxx+Rzacs8OM1BFbSNI1za09
Go40+WBDDwykkupUQtCY31aVI6WlIQlesKIYqP98PxPxqS70D8EIznFGLKV5XvzfTd6mg/eGTp29
/nqwgYDkK5h2bovRPDIqt8+CPbzYYUuZB7zxX4XV6wCtwatkWgNwvvD9LyoHHPAAjZEEC/7QwA32
NqavT3Oy0IxbN1jhpKt7yiQCpY9TlQNaAXJVZWUDT4Y0qABK82gfnkaA+zDVuNNOQP3urPWbDTbL
xFNrFby0Mb/v9NQat1AUyZEjMIz6NAGMnU+qKwi+k9t1y94NJ70QwN3Ju5H58zBcqs9o1ILfL2xF
JNXLuap25Opz6xU3O+mk+oJscXfr/uDXcNofrChb9XuEFfhFjFH9z2LUfrBHAyFxuWH2DHW46YIh
l3pno6djGdljxpNB6IvW9xO2Z806P4izJpDRIdalwhobVNmwMQ8TAog09JUeGlWAEjLRWYeg3Xw3
KuG6Kn7eHfSJ4sCk9PCXGd1fgwurPbMKwa+XOMPDMfLpYjkzu+CsuMVRjfKwLMz/fX+VgxryZzV9
YGgyYamFJPkOln2qDaomR584XWpQG/TR0/dT4QvlGSuNENhy40fCtQVTCvYY/OZ0mQv8uWgC21Ob
aN/BW4T2cGbvkP72yGyRa7t+PO9h3krJQVGu7ChsmyOHgRzbdypDBU79QDGmqnLpk/Bec5V7hnSH
BOWaO/5T/y1WDBhkKy7yrkE3iRcAKxuR1Ndd/vKq+O7fvs4sU91B27wVZ2Lm1jDHMb6lv0jADhCu
wRrt/QmWNF7NPBPn2llTr7mifllolrDFGMEKr9KEuSyvswchbLCAiQMBxxSDIzueRbLMBSsTaQ7/
FkY1fXwU3GR5fIXRW2EIn0K2qyGyiQwVcMoDdjaibJbgeY1PxlV40ZA38lLmWFfvCIuQ/LMdY9R3
hwNfLWGhlqtpRom26yQzGOPVfISMJYGD+KYqxW+cGFZ6NZXY4YUgUWZCLoC0gIUYafAOYBCSN3TB
s6DJPIF81y5uuurJUwZ/0I3Ykf2YuPCnNtze5FqWTdfZt9QGPZHHhttE9oLlG8l+foc1UOcA8iZO
GHktRCufNxcc/wYcXOaDDp0duxHzowVMihp06ukIGLc9dFZHtIBH7gvlfSYVoN/f1Vc3KZkWvzOb
2hjc6JE3MflrYhrL6eF8Xy8sIWUCQZlLBP84NqWnz19vJzdagnfz5U0o8ZwaApkEmElVYxOuvb8m
46PpXW6R6lg6tkWNUTkZol2P3o+JJB22KJNUWWB963U21fWsUf1ZYP9tpIizPC3H3s79GyUfGCLH
hhfk/zar1pFP3kbzFf3yK7L1VZyz367WmlcLjPTxAE2Yevk2p+6qhxj4fpRpccbKbCiIsFXFh1uu
msBmHSwZUvMFg+sHR3TDXnaf19Rzfor+YroTr3jR4T2ptXSwOjWI/WGnYgfNre6ItuyXJhZJJ21B
A0mfiaaAppjg81jUmD1icqHAXFdL/w8raRX91V5Rw+4Pmq9EvHtJwXf3VnKQzRq1Aetsepof0ZtI
htT8V5icYU1vjiy0/0FRNGDw+LyfdOeczOTt8B5YTBYtTWr2ihp8kFM5cZ8lu9Sthn0tewZDAjKn
o3sSh/H/dOBNVxahzDnlGIJsbptdpfYWUlkXjmEEjHKVdAceJ68jyQ7Ctrr8Y5rGA0Z6elySZoi0
G22uM26+yjikLXJmJ7Dp/eFWd5nmMwTeT0R8HurkAy+GNbjsmd845gO9jv6RXAT7lWabsbEyinsQ
33NvqYeBVzd5aeHKuy05u2uHjqbdaTHcRJuVcP09RNNpFXE03kNSTVG6BiJOcpLEseM5T83M6Izk
nPptjj4IbHPLo4U7S3VWKsf1cHM6/oNXASDPmWniWx4S40tJUbncq6kx8Ey6AO2HLDOaSGSZK4tf
VWJkLCRr0WU+NUWCZ0jrrjPWKIQczZ4xq7e80OHIDGhuW2hBMXy4vw9TlJd3bECHOdqYKN9QTU+s
vpy44P5WvwvVB87swxgYo9sp7XJ5739oB0js+1H8RAx6+DTp1lymEESFauTQ13hjkHRrL7d13GDM
lBajwAIR7bcm8IqSIfc+CvFa4ni6lG35wAjC+QJhzPvPXAppuDSdUwbg6goF7En/GxzIEpxBY850
/BDFpvQzQ3paayH2C0vvXYSrHsoZ4SgKggL7c3hv2EtKI82cSL5ytMv/4QAgN5V48QKpBza/l8Ym
SmFLJeYsm5+H3P4G+1ur03Fy2+ywkQGhZ6ctpvVfr7ur5PZSLWoUtU7WcUh6X9pqszu7VG9c48zx
kp5HhnsaJIglMc9Spj7W0dmR+/SoGy8Hr6kkMdvu8GqVRV8Sfr5gHIRRDXyD8wHng2+0CaK1mwFs
gG7tdoHHBbvBlDTtLCyyCLshoES3Gi9kOi9nvRRaMCBkj8XrPUTkZvVdtN5j4RhtS8N6x+pA3t8J
ll9iczlv85eiNR+nlOVCsL1oQ67cyc48ioU+Z47LFVePyNBTSMyRq9NMMFtBaZqGqohurgFuTxyO
ofGtrlShC43KvMWfT6t4+2RbtdTHtSNTNs6L+XDoUFwTeCJ0B9wz0hjBUZXcM1i3f6ZVpZabs7Y8
krC4BPcLejDaOmzE8tzqc/DagYloJCX6evR/BpeyD+dnG+P/ep6P/0jWDi11klcPebQDYaHw+S2G
EzNj+BxyAB245H8yfQVk2CDkU6iC/dIRAXEd/MYhkI2p9pDmGkIr8lULbgc4VeGih7rpBcOWe7Mc
kAMQ+4HiSsGIx09QDJMnxM0Gf6BQw/cNU6hH+OuKzPgqNISRb1qQbyHvDPLrK2yjsfVAo7cLeUke
DpiGo4XcSGLHwzbRsQdb7yIh4VrOmzxjpE9vR7itmZaEsKzvW0GkFc9CG7gF5ghNxI/0ngBuby9Q
AVtByv5DOhJV9R9adxH1rvg+cIjo1PGW4qGzhCP6wLC6eVgrx7O/s7GVCCKFvXrhWBTRMkPZGnpa
/Z+FdcE+iP8QvnegV0DeQjO3chQx+jK8A+DLG/TPrw3DJUmmMrE6hUt5HSrEgNlqsPdpd9Edcu46
d89KLpk2ZIPWq15AlKzDfvs8gEYmu52ouoH7K6NDIopdAUAcilR+aHG1PJrvrQ+IJNaP3WfNArBT
yci4bqHq8AfIo7dJzkDjcUZwSCwQL2OROh4MeOD4GfQYR9c4UL48byfs0RvFIA6AU+HNXw6GXSEX
QFaRD5afJ0lCTc0xb2i+BphrCi5LDff0j9TqvfNLFC7VTgiMUsQbpAYHoN/CVdLuvtxx7Me5bbQt
KmKjTaE3NORgU0iq8Hl1KImTBDmlzbDbP1EH1JBBrGgXok5DbLyMZep35TIf6jzUdGmn0JoytEL3
14UcYH0L7PwznHcL6Zx+347lDsJLY4ZcNllD/MzrwwFlp9/1xyy9DqzP/HqKjcgRN09TG5saBBBV
iBRUgATUX8qNOvkFBs8DrjqJkpW7RdEYQoWaZAjRRauiskZuw2+uWMdzKO8n5+Bc0bxvCZLq+jUJ
9NBvUY8mfXoLMLfUeewO2axvO4JiADARfMGIG5kqJooFoP5hvs4VVbNLwuxl4D4nYj5iSfS8Y5rY
/PfeJluuUWgcEm3px43RO+G0N2nXY6kolgm0XylqEp68V8XZGyIoYVhLlFO051Z545/0ynWXb3eK
vHVCRjDJuCXlqf1SjzAupVOLRiLLuhvzHEstvFCuJcHOos8Cthn1XS208YOeB8UlVSjAS2nkR7JG
ZevdcX2iWAhWfK9L1AyU+27zkQOh5yrGKNg9mKZbIRSgGiJvNyg0F9bNykWZnF0Y0apVFX74ODad
LGIPRqO+yzsHGrqIbBM0Sb9bnNoyw1VW06MPExuHyErLRgnWnQ4ch6PIQH1I2niJ5Sqhfdr1PaOz
DIZ7mqaxdkBh9Dx47D6/Jhune7/r4zALMLt/qeSJAxlM4xhKuLded6rNQZChf6/5Ygmi4OrvBxB7
7VCx9Nt7adS8Ps7ohPGUjSubXcKm2uE9HKCrY9UnEYKJPpqcjrG0EPVjcMwdnC402zTOR2TwLJMv
8POKCirgseDNysQa+b0lKwaVFal4W9HiTIDG3jQFrB00jbWZ6OREc3wBlQa17KYgQUnNrCm29T9o
hZWiMWQUkUm3Jr6VYMRq5Uwf5iwtqEIdicXCI5WU9ub0J4CMuLAEda5T6hiWLMjDnIjaHUOD61uy
EdEoWP9rG4JAqfprnk3bk4BKMlr7r3MrePDPPVz4SfXnH4Bb1HU2O41oKLr6Wc3jUz/dH99/Mqcl
u0w/5T6LO7LXLUIlm62JEbcl91Jmp/zffYT2w7bSWNRUKE4fQm5/TSx3zjULDUR8pkDT+78adtfd
VU8HQ9nti+78a0rOLUfFi2LPesf337ja590cZqWFT8RsIzZ4ixIG0fMjslqVvqXUQ8z9VQPZsLWl
QdbsDzp1LGgJHiJOUYRsES5Akvqq5jqyVfRntikOWMfjvf8qleiZYVYiZm39mLgjT07Ba7TGjAzL
daM8LqBnzXeLM7VR9KIfsjg7HiBX2HK/KJEacmxE5ZrHMGWgNiyyIFCuFrD3/lbuGGjy1FrkplBs
h09k5GIHcpjtNwDHYKkaNjwI2Lt4cIQhkjg0Jxeovj1S0YF2m0G/V57DI5jbPAi+uO+JDhhlgeL7
QTdpWZ0BOgbIwazPkP7WVtLCLzO+S15SLZGeGSBN9nWoECgMjch+JCcTgUhOG0klzYfvYpn2tCIX
VvyuEc9qe4CZ0pcNnz+1V45RhEJD+dHr/3Ia4y8SBNUUz3BUonm6+Zt9AHH2dzBZn+bZUqOvw215
ufGIYWnC2l6615hBy9dewzhJURDZD8cl0RkI689XnJGwjsm5onniOUUMLZfVaFvEYM6c4V+J4LDj
9Q94B2jD9rWPXuLI/RA4+hlf6i8lWoO7d997IqWMDY0MTjiONPFZxmIroRwb7BMpLQbufw34zh5l
X2ESr3bpBiHf/LjDqUlJQLGDl7V2gpAImyAgEt+OIXQs/CKBFqs8y6w53l5scco3wEcj+YRY+qcR
5Q4q+/X4vu3r8oVShGtDG6Bo6HyDN+2KnStCUAU3xEMgE/yPVmSX7zIWvRUT7HUCmEvj5+EOCt75
yw6ih/Tyk3wldun1fHJd4Gdx3EZrX5vJVAMAqjDDD1wo7jfwODxb5BZY8qmZk04l9yyC+4+e5kJ/
F2XKUW+Fr/rzwk+6+4SZPhU543F6pwEslbii5OPCcMNPs2mq8u8nwWDZ88lemymhva3lDTDe+nIB
IZssnvLUBDrNOlCh6tK7lNi/dJGX7FTpPg9gRH6Kq01a29uYDLnwWdoJ+MgiXbygmkzqkwwESva2
dugUi+qtNxm5T/cAjMG6p/G1pzAh/6bdH4UOWRuYcxHNSsNwOmoiQOfmAmHwjYI0nncZpkhq1ejT
+z+yvk7JNHNyJNweikHXCxgTB2EnyEw50ktykP25J5jb7xntRa+52E8V97Fh9WNS9kEq855hmfCu
y2OSJ1heXgndzSZZAJWYODvqkNpI9o89k9Cp/AUQrNQUCSrr9yDWINCjRUBdMem7CqZW3PoS3HWF
VFTeALzn5vdEk0W52mhcGKlnwEcYL4vmqkjkaUACzevKiYw5+/jE6gqHgS4D5iugV5vWGd8udh/5
/tcqG35ZwoZ0ON/sZA9bjh7YPO63vtnUqP/4fGYyI3pP6+5fMwyEOD2ni+tMRAehlGE76BLa73qu
g1zLCT0AzSlHAhI+SQ1Q7gXHr5f4FDFoWh9c41ry/rVSog1JjUw2DIJGIqSRbV+HakXL2+l0o1QB
BCImGa5t99fDh6wowhDhr9r0oaYG5L09PiAOEVwjBPtaPrLYnn3KgX2T/UDIC4pLy9wsY1B9JN6E
v8GU2vDp07+50X2PcclLYGjs+lIYKMSaN9ftHGiedKZBAOGOufbGkzoRZNcqyfuBfQwKlvFTjnSs
bA9ov7D2HW+MOobIysKt2hYQ1cGHBrqy6ZY3y5vUIZM10XlrWiV7sVgCy/GjfsBJOehDT6tEh+L4
q2rfnTJrWfo9Y+f4rUan4eFMRuByNBFAp5yydIx9dF1TiidYGunhgD31zUx/TFOLgh+4b+8rWKyY
TPwxU/Txb/RdEWz+eShTZyxcjZiCYxESE+wLfNsEpwRnM6zkHIE1zaojBPH1p/6U7DUU09WwGxso
CbV3pJ6NFwvNJAO9u8P7J3Xlvg9y8VWIw9Gw/53b8FMXTLGSM24Muz8uU9a2eJaooTuMSwhSFRwL
UISp/7AmQs4AKRRNqgPRY0tjjztkRRSapxdxKb8ID9uFVH+Xf3jIQljEuEWI9sTk5NtGmd7VDHs9
IDul8nA84pCh2BUQ3SWkLqvUHijHiA01PVoCA+rn9ZQ0J/ROw2SG7WmrqQimCMMYVJkqrg5udhkm
nFMNyhMTlHJ/jhelyK2lLxsHie5mgCHESDSlyI0feKiQum2g3RLe64EpOSztGCxWWWw+is+T6zqT
YKTyVErX5tM20s2aLmfVurzcUqw+9uJXJZgl4M60BFkZfajqm5zeUoMFkSOXzjjzgmmXPE1EQ7Nj
4GqmEq22UvHUhjtWdlt+55f86QwXVaAWyXi0tAPbPWlCa5etNkUDGYT21/06EfG4HCmfuWYihN0z
ZX8Wyo1OOgqMvvodUAlNNEPLz55CDgTPIQYiQTa+WF5sllzbFGGIqKAtKgrCozDvAE9uZvovtIGY
9zg1aorcb4H32LkfBq+NidYQP1SVlIZEXs5QO4CbXSXyMoF/nUbJXR/bCkr2VX4s1wX1j7gIBF0P
ZiDcpWjEnyC2JQahawwAKjp7OGf++zmB48UCq4+c83/HhjS4jhEefhOpNHG3FlDEFYCBveO1MsTN
feSMg+XYJZc8yT5h5hHpfaL2jEwMqxLqzKU2gC0n1Kk+xqjYlMZ6Mb0GmpglUIYDFrtrz/X2qpvO
f2pto9ZMFyuSXFgEgxUcgtAXsH4vl9wr34W6dU4Dpw4phoFNG10l99ZrQ5rKAz0nwf4laHE1yJwW
IZtkxFW12btUDp+4Khr0n9QGHsUkPouWPbutw5jBjKZEFmBojT5SbF/6nokOFFf87G6AbLS3TLdX
uMbSqg3eOlMb0RquCkVlMk6B2xqYAXzQvpFoG8HGD62EkaqkpYr4icxIiH2tCaz3Ggw9xyjgAe+9
wJsfUxCEa3c34eqhVW1vjTla/CfikT8lQnNAWoA1i0O35tyL1u38tB+4J59iVKD/LPUIY7MP07wj
M3lwrU3RBw/rmZjx0YASOveWzWJpwlvX8H9oVJOWtQT+bXdZiE7tMRgRkOJsqyODW7Q2VVIbSABF
2pLLSX5G4wPy8WrH/6lV+yGVBn7BWkAfN5L7HGDF3/lyyQrmOM64uirIOcqOMULogAdQ8sZkxNBd
pXOOYUrQ2dOmKko2BYnYxgLEWfwWgmwCI19CmcdjxiLQ4YocI8ehhA3Y+jYh2a9tcQStWDZFtKWR
I0CMyyxB22NoBjiGp7Cn6WccjW5gDh2FgF6T2sJUucFFkAZQzyy6WYbB5/if3LbfwlQR+SI7ABr9
t7G6FeQ0/R+R1baJRDdk3abJ61Dv1tDMEOtpVU+2uyAe7JDK4cwfnr/ij4oRvwJFYNfsQsd+zm5r
UAFNV9/gws8pEz0JyA/KiCp4o5F2b6diKk7hn++JNH3/HX6OblzIFFbyVVWPXQrP7G7r0gF/Sbz7
SLknvYAST1QLs4mEYzntW1VlZ3uutRJH6GG3lOXciTkHgmSNp7+bj2ack8bbf0JroP9VdKSUA1bC
A8q236JsXeuKH/fuJ2cdi+btk0+UOplcEHrFqAz9izBHMweMX/xlypgXq0mNRSlGUIC02bpIhN+b
ChiYGi5I2bxNlRi1XUUnBJtZtvrTlnsdtRQliL46vZaNH493VInvg3eouPIk1ODc11plNl7iIrDp
A5ieBaLy3+KYkPWdYh0NGlNaFHoWDnudZbcNob/8ZdXrxdzeAxY4iKxcAsWBgcCEvaDg+8OJEhzo
OQTKzlcRrGaALgi56qadMkZ4S74V5GAWye2AQi4iCeQk3HYVnuKuN1L1S3YHQMqrRH5RFdrmH/34
ZGvy7GDWjnSWvjrhzUt5sm9L21lsexhSzIXxFbjOe0o4bhOkEJsPfcIuwOzrt98VTwLGXJdAV3fu
1M65UJE3c1X3PCKHvrM4Rc+dMX7npX0+QnShgejaIiCfmKm6KR+v460b/99fgeU0kr/TIogYA43k
KIJzk+7arTtE4DL5G2pr/K9QeHihYkgIv+kiMUo43VY1xTU97rQS31tBEiUpTDswqCwYI/aUQhjW
heqp8pj1yo0HTwkQMLsvaYUNdHuLMf67JYv/vUjHWqRqM0Pe6gsFsx6Yk2zLvPeq9q5uwGq6yXMw
v9VxJSEjZRPdRE3kawrtEt3QX+nmcL0dqcDS3vlDPxVPFlQw7o7FOk2U9NKKHy45okgs5cAlXJGl
JDxpKkzcYaWC0dGb8S7OsznCBml2/BTTRKsZSZDekxoRLH76+1nzHDTzZNvOLvh74qXGz2pK2WxR
JpaofNvFEON9RkvRRSQeZGbzbbv1P9PyaJQUeFPK2q2ztOOYiYjIw1153lyXmk+f0TdBaSq5R9K/
3zLu4grSVo6KchYqHO7B/iZLSxn6jVw3gifxdBWy0SCSg47R39DVOjgZnLu7vLicGjodLZ0EfYCx
TWadXpZRg3Dr2Lhssx+sJ0wrgx6IwyjCC8NTO0oBMdy6QNLkoJYheVZFyEGiXtuJ23A5NhqErsKE
V1sJngwIm2u4nAHZVv1m1lKOO1NjfFQB/u/B8+zN4PFMg0ZBSCdSFwKAsM9G5l62/FK/h+85SFwm
aWZbTKaMS+fNsQiZHxllyrBW6Oo8wWk1oQkThTrOeAokLGoaPZjRIKRdeQ9jKseYR9TvYhYreBH4
08LTsU0ukK3FMWifv5PGZ7AOmMHB0ba2x2+y2Du3frFvXv40bhDYYtLhbJT03IxMDoR1H7//tHWA
vbmInY6JG+ZanTHCPzAdkjtFCu8djYWuRnhfj3a28ikMyZrkT8k8OvIyOenUGjbYnr4Zz2W7gz0c
q1YLZzoPCkNXgJf34SDI69DGIoO48VOMvzxQivYAqLh7xemI3DW/rzfOvaNRVMEynsnKGX9O4sdn
L2zdRUAsoBarUfrY2whyzNnvCG5jqIFiYQv45CoNAr1IIIc+V4Pgkcye675ih0FWXZ4YsapU6nN9
w2nD8N0bc2yiLI4DSauc4Gnw6F9UnIklvK0Ye1Vyzl6dIGvCWPqmTwsBb51WAw0+zLilXC0SUmyC
h+DiRzn7iEuU0hX1fVf2+coPPpeyu7yGglrxz0mZus3axKtm+mzb6pWQiNfuIZZtFvLPXZDI/x8u
TiIvDlpMjqq9awikNl74t1YMw1riKEdKs9tzCkx6eU0gmUyOlEgwoMg/zNGWnUz3jVsGTF9zSttW
LOI5BTrRDgTzPMpWJOp7r7AW4y+uiaGQ0UeiYJSeH8x3b55tV2v2hnFVa7H7HXYBgFJY9UpWEiJE
iU+oG68J/FnRcreLioCEMhSaJN8y8PfQzZix6FElgSG+TxEKHOcMJyCNDx6glDyLaGpAFMLZIi0S
t0LfPwEL0sMc+ZvLGGdHaowCQQiNgo/BfrNsTPpckC9yr527biBWcLDvuQfzYWO4EyRUrrLwNWKn
XeljK5bPvRKWBPv/bh7NHfinXrm0jHLTW/jUTbGZMEl6/tg3DOayJa2VeWc/LWAqknnuGYwrXBWe
Rh/thYZDOW9/TzZIyLPX767GnwTk1EVazPJXqAfEOI1ZqHl80NjZvEtEZs+LtIDz5dm4OEeZaPsd
Sv2rBEhJco1FNupQPXc9+CDmuX2Rmu8jTq8VGiOzCBy9CSpTd+Lv6DUQHhhAMr3/1dKgkuZPRWOT
uOs3EXPMsogV+L2OQHW5ByRAbs5fY67LCGzG9RsZmaiaDfJ7jYeYTW+eAnrfAC95NXfeCP3rcNtl
Hivn+oRg4o4Y437Y3YuvYE+exrejziB+fTzCmlV7u1TXTb7kfqZy1wkc/uXyQkYPOUgyC/faiciO
YwQWVM/Skb5m8BWPi2Kmiey4V8r7Xcw926/7JncZkdFrVlvrblI0+YnD40JU1UnEH9LlEkk9vo2I
rGEZDktUrA4VjyQeUo4XdDw49NG+RgoruiK7zYw1HC/t6nXhmUhal6PTlw1bXg3IH7twrevmjXOc
4gTG/ljmznXExsOA3Rt/Ml/ZrrvbeRKuAmZneWLSgbgGMw0LtxDC6rvSfIHZw54NcSGFmOiJkn00
AMZXCRJ8FbKJCZEZs+TkmEmZNIuhfpmN8LznMdENc1/IpGKAanV8/83o50l1VY0ioVxKmetWBZ9t
WmReE7bypPavso78HyLymFQEHgR+pCF4/0yEkv3/judJCp9EvxVWKZKfTM0sFoyUkBU9jsrw7VVb
JhmG0d4WokwSH0TxzaWUXb7u5pL6Ie0O2cR8XhqgkGmmfbHH7f7Uu++07cSiDuCKoFCpe2HtyaU2
pD6jur0yu2wZ+0UVuZs2Ie6iquC9bYFHWMHRD9+9CueUSMx3yurpSq38eqbcgXcGpFWfzEHqZpgz
ZdY3Z4z++Nilo16f4jdki6MePVBspe3TK2kBAH1XXvt/anko5DN3NdVGMmsVBiNKgS7YPseEqK0T
2z9Rvul4xbGUvrxx5OozpJabm3c5UKM9a0N2BwSEtvrpksS/NtOhBbtfgcjRNAg8EiPMomL649fs
7suggDOX8iDsTVY2hlSBEuLbAiT+G4ryrlyQWKgsD+cuX5bp1XPMEKmIm+N8Jhr4ycbndOfle+Pw
8qWtgsXKVuZGOU300jmfM55O03FCYLbmnDeWeee2AD1QMvOIE5QquXiejJDNUMz/dNQao+Zxmc6j
FvvUKad7wu41JFN5wzcc1nNVOxvjZ0WXXkiiX6jtDXwicLyvdIUX3wGq2JnDHmufDbXRNdgZFlVC
Gbrp85K6mU3+jF7zmsCok5wuhFDWbFuwa42q0w5Ew0YnHp+KKyTIIdlkjMoX1fCDrNRiXKKSlD7i
qbifbdu/bMNIhucz3GqUwQToqapfTkpOIxv0ZEcjQjUFqhN1YYelev3JDo4ktZdVIl6nBNhw2z7z
4V6uUL7IIYrt8pFckeJ5JO6H0OrFFp2k8bplsZrLSs+5dgtlmZtkjBq/wCjvA2yw8Yu1w84CtmN5
XB0R3/x4zvFEuGGSeTFSCRMFR3XDg2EHIM4r37oITjiynIxjLNJVoDnQot2PP4gDN+Sn0VuQVoYM
OJNa4wvI4znyL91JaBPZ4TXvzCha3pvoEmNf4TH/GDuXTVrHrErVD0be9JU04R+Uzq7O0Bc6wz+c
TseH8A5s1WyrlEA7PHpRFUKHtIYZwesTboIBk9F9iiUzH6sJYSSKYJKVNjws/dVaip4flfKg+F8O
qlcFq+rCtHeBR9rNViU5PSsa1ck5Bqq//Hk1VzuFV1WOmbCZHaaehmdkz5/vlW9ZlKvGbpUnr8T8
kRgkAymPy1mrVVrh8dO/0Hfv2st1Gr70npJGiVo8Ywabv1MNvg1wxsWsKw9KtGRCwFdcMy60/zEc
dwOWmq0/zMnQVuaHW+2pe3I02ioMWKjsK8/EXJLkJE+sjtUaKEaBlyRy/Zt6Ij1DK5XARdCsgkWl
pGoPG44mbs7Dt6rcQNWI4Zz30YA94g6bt0dbYQ1hNqoB/tJ5MBFJWouiWbNJDfl1IphvOPD2azbi
2cwrw+HGwLJ7J1kYbSm3SyoWTm4PgytuWjVasqg3C6m08qOqyYYcUHzal6Q+JqymN18GrOHsX868
ngn38k43QAlYcOpIE5py+3eL7jWJ8yXgw6RAJWoTnqBs8VXj97DHSpzY5dW62NlQpqHvSV6orhCE
0F7dokx+Yh5OAMxnjVU4h1LojDXnrqb2V1HlDRYi0Xd9N7H9bygw7lh+ztsViAxuBrlbPMUANLG3
eZ52d7lMcUtO3EpszRoKRRHoyOebmzXc/bKcLpbz0WPaccEvHeMaN3e3wgK1i4nsTmm2HXJbjgZo
az2SCU7rrHkWoVVUvxTRzXPqlKMpUyWHhhqUpgqKOQj1d/eE2dDRk3oxFcKsM9/2UQ3H1ehQmZce
qRGHt0dGLn3ksUm3lhX2CC9IEoyICFefRkE/yDo8pqFJHTpZgbLq+SXaidzdm8eWogUj9ZY+lo0J
fpPP+KL8FU048R4K9lgIGBE8O5n+H7lKj8RcAG8P7DC6MTV+nQmiAC0MxlXfGClbc+HqnT7wHdJX
W/a9D4Q3glsVSThXQDMPkSgtgUA6IW2WjCL3SjLOtLKILVa5kE+5JVHSUd/a7ATxJsF7qF+6rhbf
nKMLNTsmk0JNRNH7e5Y37pV4pCeJougIZ3NoRVHYwXXlih7zF2x1FvADHzH1g9HjH+QWPl1DYmcg
f8CupVQlEoH8JpbDKXEMyXSaBf2GyVbY9zw7D0mvHdUVEBjiQcTCAkx2WXAw83TxzPykolEZ0g6w
CDeA0SgRnK/7otfXNJY04H7qfUBk2D+QZ4u1rfxMG1NH9AbsPzO/I6bUG9SO/Lhsfe9EICKWCorc
KWr6ZQr98RYST9Fy6Fto7xltsIUlSh17zQ6VsJ7KIL0CKb1uHEmAAOzZbkd7rSAy5lTuCZbBNUhK
gwCwwQvthkPja5l+BzTbqtcNsLjXHiZ59Xe0W7GyLi+s69Dwmvor+x+OsYcSbodkEJOB2GHmia2N
D3ZCdIo0diOIHf/+VK3dKS3EBGkD8a0DXiIVfEa+8ALHDHFSbF2qEWEr9nhu+5IV1n4zcp8vkrwJ
dU0JjFWGhtcQJoBiUjTBfOBOyCtJmVHMMre9TKRvquIBqylXmiKRlic9I4/XaQJTH58ro0cFKfIZ
lG13bZnnCFnQJaFHPn6L4TWVCv537tR9mRsZ70zA1PzEwDSpO6j6S8qQEw5HZZRGSWxJMwP7hmqN
ykFY32e3aCMgQ1eqQ/lgqb8vTqA9lJIqxRpViggKYfrlH8AF0V4e5Sn6OgTQKqVZFzoKVOnXDUM3
QjToYXEVOwji+Zu5IaY/AJ3MJ3znkWvtbtIkJxEOydA91JJob+/v9Ze1bV2DETugNmFftSbGpKZe
od1JIIFSsgtuGnRdmIqzwp/GPbgWIntwp+JepPNqL5C0tewJY2OqnYCIzzV7PBZUyZD8o8sfUXvi
F1Jsr8v/ebhqBWXG3UsUemCKt222Fk58R/9Q+PA62ONbOdVeEn5gwGxv0swKnxfgT8Q9wrtAKdHt
JiRWifXNywuZuRMlC7R88ZtZY3RUDL23nNldZhCrp/0Djo8xr+9NRnxk3LnG0pzDRDaN1UE09Cw4
CY4gFmxB7m8vaCvHuYxC9EJb+95A2cGoqjmXtO/CuGk09V1vDIkDeeAPbX+1blD1JF1K8fMW70qv
Cx+ey7pVJiGtO4tENI82dVjRp2m9R/qnRhJCs6oZ+y+VBAdF1FgvI+imE6CTw4PDG6UwiOmS5TF7
IvCC0DKHLc7A/XUdDFkDXQpaXPnR+2C/YdzBNeLhSGcNBGOdtzGzvd2n+PboXidWqhFj88j8OFgr
9OB1MkDwHS/+h3WngojvUg45vg+ZgEP2xXuzojFvpTLzcmOE2cfo9WMqpUBwaRt30C5/gZ3qfK09
Zjz3AmBUf9jyZLQLB2tUdToH2Atim748Smvun/oW43QACUELUZ37PMvhWGLCnYhJ2PV7mbNsmt49
wekSz8I2tjKOiouwIjSJWYntI4m+gA998jTAfK+zCb/wSVRa5IbmxCQRpQl0KDgNI5opNiM704LH
s1HLEVnOEG4n9jO2ZY6RLebXDRs2gMkbXw+DsQLowcmzl9yr36YuNrnTBp5dq60FKupnx7Zf7WNq
CCk30BuwKZhYW32mDlzshYvf+CAxiWIKoXBF0cKVqzVlnA8pWeJs8Ppz4t8dL+LUs0jX1oCw2IJP
CdNpr/11mmunlp9g0VqSIS09/e3ZpOl6AgVB/8uItHjn3tjugSk3hWHaC4bjEOuwTOgHSwZlcbRJ
+M5NmzBADR+S2mNOZf+qaAS72dgO47WZ+4StTekB8IP/JibuPpc/GXGdSGBSZcPScgtUgkogbcOO
87Uv3C4y6DVUjX26OitXx8lAuPy9UUvxEzNI2uYU1GEe/DrD7ACrKR/kwHI4kEECMczshC9Iwv7g
1kNm4UOf6nd4dyZ+28rH5h8MGspG4kz7YQU294Ro+ROP4Oqw6ianqZNVXrkCU2sgJp0P10oyuKRa
eUKSgUDS6yG/SCdh+vhmOeg2UsmY+s42fWh6n3OyT+Ruo9jXYXXv0vNyyYmldVnnGJo90pmJYCRH
ns+MVHVJ4mkn0s3e+BDi5OBBV0DHd/lVwz2nuNVEpz9NIdRMZrrDPH5dkZfY5JGFA9rQFS53xeit
VEnNfN1P4qimKnwgCmY0xYw2Z7nE6Ut9pXydSoqfl9SfsiLl9xIvAqGipaojolfX5tokdZOujHtZ
/O+YWX7AdA+6fSvYFaMmk4NxONqxcc79wU1RPl0WVnPCVaSG5ObuRiWYsmFEV1qW1N3FOtpcff7j
Qu7JQZ7yP4n8KW4jdhzfvFEBgFJ5BRjKkdsx0fBxRZrhOsTsvdGB534k4RsqTokv/Vu/oSsh4jMk
3zvELWQti/RsSpOzIuyYKdcyeWZwpk7RCE0n+3JlTH1uXGo2noXRQwzvvv9dtY3eLxoDBxdlsTZo
5v4+TVuMucHTGmMJuiP6PSIJmKBCQ929c3MtSJx4qDOETYBrvQy7NTwZounbxEn8sa8KX9iIw0yF
eEPaxYntLX8f+NT8uTila+wG8jISzA68iwt7J8OQcMJYLAVf6u5JTGjLfauGNi9q3vMYJlT7RsDs
sujO3xVRoKO09Rc6MyIJz0BEHjyap/mZQ2VYmZAbYchGWg6buWfgTF3cu0SM+8WMUPSvoe3w9xeC
uWhljFlpLhfjEdxPQDmDM/fRjGJV1UEaX2qtKetlqHUQ2Q0kS9SqYzVu4mQZUK5zI+CdBQ1c4UzE
2Xw+VDXwrqqdMxDyBfDYQ3DMMkJFj/zRcBkKGfHDv2g/rD8/ck7KIH9Unf+CuvxOYerKdAHOLjt9
Jha4P/1l4LHvCglw4g5Xgh7Xk6KGH2e1afCDu4nESv2uyt9DqkIg/BWQm2PMammDT9s0GJoipmqR
2+jH8nC8sNobLm5VW2A1rkKT8k0F/FMOyq30vno+Noo73qCUMucJqxOEH2IeS0z7rDessBURe5mE
4wNZ+EwpHHFkWFh/q39hU8OUQgpzvaKLD6f8x+NinpGV5NzcAG/M39k6SvvhDUEyJvXXEpB+JBNX
7wo8WgsBJ7hfdOAFSkPo+p3oKb5FJLGzsUh5mdjOf+wO9TbNDGfLhWfrCwenxLr4UnnXcOySnKx/
oudJW2jB3MDkpl82E2qqSnwLRJa/TDcxJ7VtkOypukaMnWuQQP1bb7yfMySmfxYDyK26D6w3FwHa
FXHKtRzF+BxsSOqTDlwNbl9bo7KuWwLI7l3r2mbWuMK7SvQcemEJikFccdwlAcm0ZM08TXyiPJqo
6GKNY6ivWzJK+BqXGwHJLnCp7YOx/LF36r+0tgL8QYswVSfQdoMcHNxr3HhNKECdbXTaQG73aF1E
x9yC+WdkmZJLOcMu84wpi1PqGJF6XAvFLNQxYbxTRHqeIfUkimBem/f8pudg6EyOGk4sR3PjVDpO
EK0T1zv46N9VNCHEDrYpuDcNmOThE4d3TRKHnV7sWI6FOtiU7fKe6MU+HmtshQE8e/SZigIcyO/Z
YvdOSpiIxqDsHl/fFN78qvqbpe6i4WF5yZYwy/oL4kLW+DB6gcQTmwiRqce2sMkh/8VCh3BsNPRw
0zHTS8aEvIJAC1rksb8MlZ6EdPqIqFPOwJ9bBas/dSCjLa/Afbj5a4x9BODYgRxPOmugOa/OM3j4
Bfg/XvFm8ALR6nuSS/eiWgG3cz6on8b4iHPfxZK92bR/0V/jPDmsr9J654Eq0M02O7jMyQotGROq
Gp7ZjKFHMt/X74qSiqDC8CUBZxXgemPyrTKx5V6ruvOExw9FO+OAPDZ1yiPk4NMy+v6+IqOPGBp5
yoroNJknQHsg9VcqF2SrIhWk6By9FoUmwiA5LkU34/BfqAsW6nxME/7gyj7hzyoSr560ojbXIGYr
U3kZGhwYdWQ90wRl78ItUC9y0J3XTvB2qn+YcnINnzNLOeWCva+5v61PBY5+5g2yhy4Fi2PpKglG
P5k/K1M7sXs2Exq7WgJVdsXYtX/0hZFXNwucJ0xP9XWixW/W+ZedjtWbIpU1ElWzHeKxcRzWkmxY
Wf4LWmLGiTp+4etKmBWN1HZfbqvxTQGItRdk4SS2Bv0jIYacm7Edbij5LEv3E/eBKFzoMUKD86Ys
ZaS5q1dElp/MoqJi6jr/rT20GRAPqg7GpU5tHJFsmanZNED1RRGXulHMAaniZGomEW2b/H9tnOv8
SN4C43p66NQpuJAZewV8BankoAQuA965lF/M5cXCDwPt5p/xX5+nF86v0raa8bJERUqtuDHDBMLt
NP1MtE4Ac2tb9B6N5GJH+iV/6/+7EHT2DACJHDDWJp0HGoQFFUMdaa9NpDdZuDDHu4ewUUqbRENr
GJ2d0MRYl/sR5vIBpY8VaN4IZVa8XOUTNNt7IR22TNbjHBBueJdl+45Svz2WrngVSdRTBFHIhr4S
7m1FcqpFJuyu3TxsulTNq8ijrD++4XFqOWe6xIhl8KtPj+QRGwwXTLSanmKL9mSdzUR3bkamf3kd
hBZf4B9x2IIvOeHABqlKdzIsUK5Dq6DaSePfqoN1rIjUFSdbZKQZvs2+U9lSLyx0m3utjbQTnNmM
YGrDcRI3KPt02dJSd38khFYF8qNxzF90H71LUsRiXbCVm5Rk6ESGaVHPWLzeLT8B7EqC6rhF/pUF
SoCCOwCCfgepaIqyTQ/sWmHRCTsIAkqZPO0H0nM7PyYWYdRXFxvtQEwCYssEs/9DmSc7UbcOvQdy
ipJs1OqwL0WfHSb6len8labcL+ElKKCdbLMvAGj/71NXaKVNIGl5XDHtHV7bjFi90qUmseCJFigk
TB9UiogTkBNNA3TjopdhYhHqSQpKgKsd7LRIl+n/kJHY4D5dLWajtsmMmX0/kvcb9uUoU4UbCPv2
aOWoA54eHTX5udy2aX2d73g1Z52vRabvYlxlCCcGnOYzDW+pkWogG0hB6xYsCDW5UVnbjoTNgrHl
FeABDzgMEo0gJQnXPPARiAZXLPlLnLY8+9jBbzSkuX8YW8Pv4ifz78vKcK3/qlgx8wMv8BJr6Nx/
hy2/TAfJ7KAM1kTkAo7JhxMl69fr5t2nAy3AMd0lnLLY3AggkPTKKWZN7Zya1l4ZNt+98KNt8WuW
1QTfkbvfgX2VXRKckS19dbDXZ6KRIS4gKDsZbC9abHOIb3PJKCVEc856CyDqSRgcERd4gHoBltoi
esdFhXqnU2gZol6a7+JThH3N+icEih5CN6QI/hBScs+W8twRGQNzWtMMWCcv5PE34TMf8D8rw27t
KRI9agr2Wrdy9QTMcbM7SLelTcxtMyl7zATa5bmWcaD1XplWSp0M5Vd4W/KNLNNKsfeqeNu6OOsm
VZcE+yxG0ZRV9pZp+LA+O9n31I5LrDxPppKE9oc6Qm+DtQdEVFAjjAd56hGa/UmiOwkZKB/CRwsQ
AdtOyBSEhd2wqQNTBiciIsT+SeB8PcwiykZwmLZqJciKIzq7A1Wb6mZSI9w865vFUAKMiuAMxH/i
JgJ+/EDgbA/81idpeyQgyCMWkWoVh52ebpL04yL8YBXPdPqCcvhoYwfOA+dN9yRxbrqusf9xHRFb
HiOUNWQ8hAmSVYQyTgxURUG5LCPVW2CDbDZEaeDodOTHzu+ER7X29qzxZNXqZEGFx3Ea/CdEiqat
pFKQMmhD1hXBzP9oms86dnq4n49m4yc63fWzO5o0hogZLo2Dl247ohnKpWk3RTRiP57qUY7Q4qUP
/LmkLm1NzNTBi9i6pweMKmUrK36rCL3QToqxIutxdpS2w9A1Qpmbqz1jNmXsCF3ojt4e9XS2NBL6
doUeLfuM8h0FSc6T4XEFRTz3zRS6a8u+UHOTzNjTAq/MzbWPJzl68dft8lSbaYevypljN8mlVSyl
9bpA83F9Ff+kppVEhnt/5opy3xrLji2Jp7fiLJvMEBXH09U3pMGJLUyrhmHrkwnAuaiLyj0ASI7p
CZw6IKM3aSR1cwHUTGdLACHf3D9Xgv3yKIvqdeHM2VCQ0SHs0t5kFlwia/MrICYenI9BajXa+rDn
WzRMZWQnQ4bxLKQ3qKUnqxyfs3cTe/UcoTkpJ5cVxIFMp2/bk/RsGEdBMaafk/4S7m3tHunm8Gna
wkxpv86ZRJY8NeU5cHVPvB5P5aGk2b+kbE6Q3hucRvC8x4OUdN5d9co71+Tix/TQzA7L0+mGlucT
rP2qpA6Tp2ohSI3mQkUTE99ZiVpX4g5Z4gCgOKvZu+sEtRZE7h4U1aPP0GxsVx9BVvS4N8wl4btY
r0ykrJmIyy/7b4m4QxYR52I+fpWfegRQ8pjp8gaIy0bdXtJotSdE5dJNIaZ+T75KKu+GhRpRQ2r6
+ciAmbqRyQcSKsC54lCqdF2anXvvXzhTavWHzjzTlMSlLxY+BicFXx8abTSGJ8SspC5kfQqeGspV
B6tYoao+Mab+dxHZ/FX9RUv1vgqaqRpxtSBl4kCbhuBYuQVmvv4ktIvH8jZEj0O5mAsxp4r2emT3
7D7PnOsyNDyCXf+wfC0AOjFgVSmVE3PI9Re4+dt94BdUutf52AoJTelDRiwkkS0pZBOJTPY0im8G
+6ZeZZZG1rhByaG54oQB44T3U0T5xBRkRtfF7CpZjarjDJjtl/aMtDsfzh3NCpSNjD3kjjjHgprJ
WBTbzaKSQgs3WjSPoIQ53waygZyH/B5e1IMPewNys4wZhecUUCyaAVqehTERaVWd6g36CwZwkJDp
/SJ3a8StEijujZVaVmU2iPsC4w2kGkRJrXlJtXi4An06YVU3eVsdYFy2hxbPzuaiRAHRS6zL2rQg
0na2vHsIZWZdibtp8xo2EzrMv/3uUyamhLcnAU0mW5T362ANok6G0E9ExvBSNdA+L6MOuCgvs94c
KeJPxEIoorZeDpZIBmi4xadc6x4YnuUNM+gvF+Z++mvqGluJyYBZ/kvuO88IdYTy2/MImRJ9WetB
v/hIHzq2sFBXYItKmSl0h65YD1QTrBWh33iblxm3yYzMDDzQYFS1DE0KqFekeMGKagzczHJT3gOa
DtHyshRbZHfuJxXBamx0QcWPVsaM6lLIZ7S1+lkFCn45TQdZrV9aXT4+F6l+da3oBQgQ8CbPfpPG
s0LEySuUlSTNVupLMg0zqQMa5QtpgvI9uYsV3k3y2CCbNwRMC3WjAHPs5SwcOA026HzdS3pgTrMS
a+s+OEnec5WikJQEQ0XLc4hkjtHe3IUJrfk5a/O/MexjrCVUQstEuzi9/q1lpFBazgXhaSlQGyoT
E+8/JAhUFVnXGAXC3QQAJHz82mgY9sAZpTViaSyB7KaHKMwwE+pwzANznRKekgy7wFu/iG2GkAjo
OdFj5Qe6Xpkz4Jl/CLuXYXmlMNqT1k6lpa8n8y0SVanbNBdc/iLSizB16GXbJ+BGnD+XtSRkUll9
X68zlG9LYKelbG5pORUZ3S/+ye+O6GQY7f7CtHEantXDhS6PoyX/d03DzGXXCwfU69PkY/XF/rCa
az1PM0+CtHA0H8zZBRA1IX5ik8nRm4MYf+HSFGaBBaFNcPEKGEJbfVV9i4qi9gH617jn3CmVACmo
HuBf6Y4loHf0dWgT/dbNmeowGeJ4pX7ct3E/zKxKqhJt+Ey7PVWIzgxrGugRgw/qzWaTmI52L/iM
xagZxsGx9Ijtf+sl+peIEQOeskVAkjnNsVIe0dEod0z0XtdHvEkyfknSgsDP3NkufMjwlNwpwNw8
ryOPp8dEt8yRXXAZSKeVO606jaO7VdoAISmLLgtrRuatAvS6Cv+Y6VZ257ia/UHJL+TebnfTUsct
d+ILgxuPLd84wyiyuhk9QPmP9W6iDp8KI97u6/v4CsCk+9Im6rqXVKq8AAYsQujK3ymdRW+s/wrq
6EVolB00ahvRczXFF3B7r5CfM+00xGAXKeYKENZeeoRQcIa3LBmMtyV2b8fo2xikxnPZFFk4kop3
ihlbhw8SLMZezyU6I2sSck+Ne6K+azLU3gNYtbLSMy868w8eKHOZctA8ZONhwhcjfQlbhJFPayov
9pla8Ahe94zpoXXimgQ/xsar84LRjuojJxOHUhhj7dpgFuf1t6xjrEOpfCLSSqgH1ChzbNcbAouv
46IUNQG+ARIMSbinZ4hrumIq/Rg8kgVO1uGBQuXWvJJj9QH7nHiVLR9WGiJj7/7s1Hqsi6RSoxqf
MLt72kgHukgoBdJBFwfnqvDoQ/TG2wTBOgfYk67T++WrvlYMZYjO+vi5rYtnj8Hm7dNkGwSftJtf
rBjww+tHQ8jkD8pxpqcnaQTYudDHHeWxWwOdQCCntL5FbYqyCgT4dcywjQ+bt3CYa3A8sQMU1IBk
pmmCDOsxRZ1jSMmFyOWW7qQa+lbJL3ar0No4rf+Xm8DrxOsJgymsGfpMIrDrKBvY9Dl0bd7jdjQV
zzZr5qCy5kSgdnwy31kRTzrDDvurtCoDBk+yQdVmGuufX60UAOefHrP1BHIpJqsVAh6kIQom+S5c
xrQf2sS102ixgQw81HcC2vUXWS52L0QJsGLGs5JGodq39knWzO842ZveeJdJOMKKhUi/Zt9sOB4w
ha4I2SKLveR/nf9VFEC+cmUn/SQ2FnIAmGudgFqqb/WR6sDRQuqK/rYL7N9mWjHTfZ+G5zEyB7k8
iatUDYMFoNZPj8isvoAXBYCsIi0N/g5F42MwM0ooMiASVty8p2lRcOtwGngdD7JB05/YsRbvZfYf
6Bazyl7SK0ZmMkLyVbYeD7W/BtKaOkameuvijNDWYg1/ayE4Ai6aPRmnOOjiKDp/R9EZvX6BWGUm
P9pVxBCrKMPMxigkjnQhbGry5ysB8EiBURawEEweYV0ULp81l8HaE9WlGMtrCDjKvUv8ptrStfWC
ah6VCqEIXT9cGEZLI66qwsl9sRg9TiwB6PsPO1sWXWTfddU56ZvmAEbfGCzP3gB3GP7kVzpUKQMc
V9PTCzE3sAfAntmCM4VcomsOW6zrU4VUumKnMX1Nn6xENXbrmHoZiOYy+5X7QES5ubGjL/oGJsSB
YetQ9gQQQ2vKDUIPIo5IhS8oELSUp/qqvh+D3ZTRoGoMhOkrQXuCMxc+/hTj4qIh8nP3OAtuvAbX
ZaHDZeBlGCLhZABesNT8wN1cORMFE6D60x206qDvpoRDzcO5SIBJ31E5huo1pplqYkvKMig0kTik
49lUFwjVVjV/npX4SkHpyduCtVgiA/VGmRHVRQPhoVFomSie3cwUDTkK6/InQKRyJE9z/5BjOQXH
cGAaoEv2gs0bjMNLoRb+n89TlX02QuRQmSv73vgeW/ZllWpqAyIilaVcAI5oL6hVwDXQ6/1EO63D
ccYDZ4Av4sSAkw5JkzWMC/2YtuoIAi60JT4hPL4ZGwK8h3OpNC0HS2DaNZKGrFoNyd1mjoGoM/Zk
mAKcwwFx0zXg/19wCXkTnKfgLI9MRntpNQ0YEkI3l1kkJOFR+I0IdIkLHmwqrreQ06h61m0F568j
UE6H0tpCHEjnNtI0sVtHUkLbtwGqdHH4p3dGTTD1ayLB7KYEOcsU2K58DtmyWG1F1v7UOsF06ls9
I55IitDIEVO1gxJRr1ICF9I3nfAyzFi6ZwogRIOjJSDShTqTrK2eCWjvGwY2RJQiX+GnHRcNqYwt
f1t7oPxw6n2wgjVTljvGZNcG8+28g7qpQAJ33xm+FbS9GV9CrvKxzLjdytNTGUSHsD3ouOtmFgZP
zV0/CwnEdNAuxx4sdAdyUPV/Sca90u06OdO0FNANW9tVee9oi1X6+8W5dRTL5OqPgCYK3algIAn2
3VN5rXVG2HnnVOkXugscvH/fFeqmyNobxe8MRhB+W02QFhy0sL4K420TmmG3n/q7zNuiFXxlKe0I
a38+Vfe8rAhalYW5R12hia7vdqiEJJrxgtfCZSQRMYTkgGpmtQyr+7sipQ8EocG/a4H5cONoUNCU
p/1EQEJ/UWm9E190r74kXo0XYMrh8MN2EJgo7POQ30PCmLKN9KKQt5h8r5wA6RGqJrixRguHSSVk
ENnd3q6M2jbbPOQmVbeanIpWWqDjb2Ni3/WIG2UQ+3WbViWBWkm+Nbs6wc29mDT80PRe4m6jcsY/
veflTdDf9qhqca40lkZTdefUgttl+ohCefCdWYEPfdRRlxcsHdemAI7xizyt8Xv6QUMz8PRocjBf
sXUUT0kDQ4Mm5wyM+sXzJJhGK4c+4p5dA3evu15VDPvJ0Oj9iLUWz/xIXyn3wEOuKT3cWhWo21rf
ErWf2KWkl8Vpn9VfaDD8+JWHDlJ3tyzF4QcbG4njFBcSDonwjPzIlrPnwoSRaXdmGUFfJrXgBK9Z
ZUBiPPqqwERHaSGuuqOk3Fn52EMzuD8K2NxdRWhd+ZqbVNSlaCLYIaCBtkzuwkwI47QHp/USiLXn
1ed2fkNvREh5fqXh+ATzQqEctLZa0nYMZ7Mo/3NpGZe1H39uDDvjl9dK3LartXjQzySlz4NGVdyI
krMWxs4rwBGiL8GAJl72kvss2QWgy/zW6GzMkTO/pi/mcg7j4d2dTExipTJcKbQpQBH4zsoLSFbi
BJNUgYign/0UPeFrDrzSU0UGjYP5/pZgVspzXLY0q4sAwArxrw7hMpuHqpi9E1Gqqk4tv46wpqId
gag6RPycWMCRde59PBhpPFrCmVGhrR7qqHnFG7vgm2Ce+4QY6G6qUJ9tzO8F+8xnFDYTcPmMocCZ
l966ojxyAL4iQfVzY1+qmFtKdn1nFB4GwokshILMBaGVO6L5Zs8245xpOxqv82e8nAwpxoqmk5z0
0pelV8Is16gF9TDgvSTj1Zs3CPVVn7T3maMTw+FJUQAtoZuaZAW1wNB3Cr5jRX4PzbQT3sV9II0Y
hfaXviYwb0eCngamg7NoCrHbvuqBfhg0WlvwARRhhVnsB3Ij4RmCr4UOmyIbJQl6Yla2PtNme8Dj
AJItAf79l6I9VTP9pg1dPcEBy0hdRTpfDLPJN3Rbtj04YP3J2OcShSHvHamUlRQ6cBpkl4YZRmS0
pQuUEQLh/zFXjVOfvQ12xHPQ9lW0vuCD5GlYP5HDM3bXEseKETZOaHrKjBgzQavmSJr97TJXpZOm
kO5vnhpN8v9vCivk4KmGDebfWa11+nWuKVXpFW7XBcKPvm7rMcDV7PUHYLnf6uS3tpAzve1TDP+N
ndBSA9juiRUZ/cdnzYMgNsXID5Y9vBmweGFTtwd58CdJqM4CLyhEsggxh0Qow9kuuKMHME8CJ4Qu
j53NZssafipG83B+oeh0mIyuQjmYlq7orL6aJ6I6U292FBrZaYwtEwOXgrSLkbSaTZLU6yZCOLJo
TktJyCDkV5zW/i0Dm6L3P2kPBN7Qul7MOVBQKilFEVP94uXJCaRLM4HJWbYViQTisGmMLmwhFnpQ
LUDwREsSCE6MRHMO45Lt+hz6O1oflK3G13pXJn5LI45wLQkFo/boNLBsJ5NjKIk38tFNQSQ1dE51
kMirG+Hpt1DiCB+Axd9xKz40rwvuQGciwmlDjhlX/ULoj73W+J3OLscLa3KEcXYNXw9jujMwlGWG
CuAtDA7W9ktwgCDiVBHm1KncW4ttre1GGUxYlgTw+YcCDwy+WrJq/D+MqPwoOGHgZwDA9WZ960W4
aA4caM0Uf46HHnTgWnQqyKMAt+lH40XISXuzl+TQ8B6+hR8d0Z0TGOlLryY3UWRpqcQZM2HNJh9U
hcV+tChjqwwVTDaDZFywjI7NjCEZpjX+zrph7ykfk1gSd4SBQ5/lP3/Dkw25nrd8tXtab+Dz3ew8
xaeRNvUKxy7KsEJUkqddURn70K0lnlX5BHHVnlmAWU6SBdtGYLTHDdO6+iEezDQSH4webmadIl+q
bOstZI4bAu7GARamMqVqzO95hz/k0DUWasxMRDsY+X+JeUyuHJr1S0hy8BinaFEfjTVDiY09OnhT
xPJ+/y/kd77dSv0aQNIdWZuKP6aFcmgKj4dlZ/xz3DZRIiuzFNaQpTuIB51nZR1G2odKTcmEzErh
BtR+GeINOOAWcUV8MBSF8M+pbO8qm7qIFxmvw9t14Vt9WxyZxCjjU1zSTnfN6MtI2QHZ6RUQ44i9
Y5nNLWT3bVziFmPpWOU5dPyQfOXjaZbxby7sGbjRRjVwDQiPK7CXihTnhYOvZ+FacI636wN72xHc
Q7aIYaOsylLgVGM8j0QpTmtaYQTpTlGtISzph3Rr8DwrcbaKbHauDwhHeZHVaGJOpYHK1TVrJOar
m0Mf33ygKB9h3kYDPulr50GO7wqaks4aPr5BNJW4gh+0LcrGV8/P45DIEdyzQROPxkgJKfLIIvfT
+oykI9tHP/brJdivtCGuaiJkdhOImmLpQgFSxAkG89ap/dijDe/Nk9yfuKG9hoYNQeA+NmtEAOxp
7vtUFaUsGSk50VL5uOM0cDGj0jffPH0Xj55o5EVdPd4qv4HHVJvF3aOy75qVqrAE21bQExNvNYY+
4Jjej4DTMmKx+K92e10MHS7uU8ab1cBT/6hsbLtFbS9huWalJb6SuNyJkYWnovx1T9gmidAYh5Wn
+I4hG+6d/YALMFZaQfG0YGVhkybfGfc4fvG1BuALRQRCe+yiVGmgpi2xLw6RiU6lV1HlryJbxffG
n+3I4GJIvqp8IHuhE1GLOqz+LTNF9vEJN7wCkFF6LE0vVsdKnBmqCm5TXAFwcDW/vvjVvcPhlXqY
Bj9sfxKS41m/7pc2D2WuIBCuGv92RpPY/3ZNDQ3s+t9vnKgM/mxSzIMb7arR21KGzIfBWaKPJ4++
0X5w67hzn5cf1VGVqgsUNj6LwExK4j6Vx7Sd00gyGejmlfy9U3rp3pFMQcmZ0wTjbRzjQk+MwF1v
8Ll5idX0RegMVsXICVCbkqhG58qF5WzNuow5hVLZFcoZs/3rQ21sIwjKWZ16ILdmiuSQUQwoR0MW
SAHEz98zf4A6MViHF34CY4zGdWJfFtTxLx9r1zMzqK4sBws2hXbtoNMDp73taWf9MBy/N1fg1xGq
OmwxKGELFbphrjazBkfmsdFFA6KKZvg80Zj2dRKaS5AvkzPZfDoB1XCL6auAr9rHWXiXMfxcyKpr
4qF86ECD46m4tpfnT+gYOiVkXTBAs7QeCenqVJK2ytKBOU6oVCQpVrFf0EbK+MX9FbhE00HoynNZ
+gZQaw9rwDiCy28TlzgR7ADpk5uemNVrqWNAYkyuzgmToSYnR40iIQwgCVuxMg1shf6MK1b0vH4m
buSJ/0oMhlB/fTPKk1ECNIunw52QZGleuJTxt2HK/CA4CGcG4BTBOQxnlXBjYf3Qekvage4P8OUt
wndOT8fSmbVIi8PG2a426Wn3u0YAmzw0Ds7fkD9ETn9TDw/tKeo5gv1gs2sromUwJDw8JDjYwzJb
7zel1LkVM2ZcMt6wGfOUusbPhwr2ZQ4dy1ny2AeHAEIhNemlCPtBJqYY1XmZIA+N37AlyLubaW1S
4rhV9yBJAmlJ4+f2i405ZXFk3HZccVAYGstAwLrKFmrvSHSYuvjYJXhXCfWUk7NS5NsuAAQIxvuu
EJkMGGbnNQg1iX/gtCvlskZFRrgCZhiEc4wcEx1e0wd4QkjrCVQfWXxMXfjRq6apuZi8n7+gKaDs
N3PYMImk6wroKZhDcCess9o+TEkGty/KNvuuxhT5c/HJ2n8lkp+mJEA2BswwoUWmKTPEMZSJSJtZ
BFt/LYvaAJ6K0oGM9KIfprFNuJmi0u5zi3ZRoGCiyVp0lbFH/CUwPtWWGnQAwD5VZLlKFlHe478A
omBX9FXt2GWAgpN2RxKPzvf+elNUl9M1p+NAWrrGpBN1nAeKkbgt5iyPajNZsskBv+WSH0dIikBd
VfIz8pb1kfjYdGrLh7YV+EAkNHlxcdiNi0gSPRs9GUZwEivTvNdAYAEVAR3ujO1aBdKFljBsQAVk
u3wrxfyMF5MaKs4B6jQ8YXgtoZhU0/FnEZYfUP3AGB66IzADgSjV5947fqeAcUU+GkEfosr5Kx5Y
+JQCWAl3phuWqlKXuIlEIc9k2u7XCIEi/h47Ya4B+czQ8Py1J5a3dvcGFuiIX7ACR6MmssII2g7E
657dbJC3rcTa8JGiLcjeJQlTh1/CehWww4hP+ngzhSFpbBwa0ioSq+NNl1IDfs/M6Yc3D/zuXO4Q
wC9H9FQpT9tht2GYNMNq92Fz7meBUQWLFNyiV5SRI7DHZV+Eh9W6vt88HNWEcE7oOi8eUGNt7tZm
atvCtzn1egv5u02lJJb1crUC3/9Kg8tcEVOwaNjLpt/ErB1/mAAanEfqIBSv701WupvMyPq12BVB
HAusNeSSsg7AG7ebnp53FlPVzHJbLGnQDLy4LrTVDsRKARykNSvcl0OY063X0KeausheGMaRPM/g
+4QNZZ91X+Q76MuTBYfXMZ6JJj93HuL4fCiKjhSgRruQ49h39pii5davcqSc2QL85Ew3j76nC03W
a8tOoowImJh/ZWU48LpDeMuXG5wk5H4Q65EjkNP9kLHILaY3MUPnnwAksKNQlp4C1YGuyZuuz4vg
Syh9HHZtxAxi2kEFem+579y/4CbLkn7mJENSW0H5X/JTkix4oz/56uUjmmIjYZ2/dQLmrrdvlNq6
EZbrnuW72yGdSIHiGe7bR9F3GKFxiFDpykWxK0XaZgJLFWSD5hygbtMjMkIPkWRATohO9ViBhJBf
n5aU+/biMgMKy2kxTqgqVTCAgjsOYczcejsFMhceeOZVThfcRDhsdIVVLvnYtLOKt9b+wOR3CiUz
VnT8GhbySv1Ih0Ptn4jtVhrB/uITDebr+MbjsYa7WW0UmmTmC3Rzui82fOqYwhvUy14PXNvjOpcl
CmaituEeuBHjPUi0yxqD+bXSwbQBU+NEgZ/JiT+WWUBUfPTQLXa4fG4rS6FU9f+kAW7U1CD/Ehu+
CAidiTZcDEvQ39AejB26m3Hzb+4cX3ZPivCXQwpwEsxhniumOirUOvPgZRJpn+Lvma0vwl/ufyVA
0kU2AeoNTbUS1FvAkuLWjTbZWTQMFSYt9UfjwPgmSXrMLP+ag3g2qsW5nP7/IP/QWgPq27CEhH/s
oH2f9Xi84S4hdjpFyVnRX5ME279Iwq+K8Zf931rZuf7YfSdzRobk8L1UOwgiFPYrbvP3hoNecu3K
6itz7/NExmOTVAVsGxyCgE7pGnJmY9iGazM9S8PBCjeYK9p9BPSzkJ1Nd3dyrNpzoV0m74xOyfuj
kvUiysKA9OlifHKoMkB2/7uq318vB3EkV4p2uoHuBwkOk6JN02KXCvqEMQZmKXt8e1EoYhRER9DP
kzTQizoELJChuKNEXPZVurGVjPFASu69iBDHxxk5q58hq/Ve9greFU8o0arqDv+/zYSwNhaXgfV8
z73feC8at8zjIied11KMGrpBGf3deEiKba44nYnby/p5mTz6LjGE09ZRDvEan8Qp1IN24Avl+38S
REoePnaRZSJG81ZehkrzC4qSbehdSP4iWVWvvKKbYWMdFn/NdK6JOhyaWx1eCPwr2NHbcZgCspio
y0vxXBsWcw2C5OxOlN3QSXeBGlNVLh4h/N0MQxCHlAMOwFFgNhebtOBcKKXCBdM5iIEStEQRoeWV
Ex4Ege0fF8j+/NKZD0zZBwG3U0qjB3lhlTE5SjecYqD4XcarbSoE9BPN/JEMK8gsN3iYRG+sbqXq
YwdiV7RcXVCMkrWAuHpjv+SQgIWXEz3ErVOG4glaNeMjw6ODchejU+tkVthT4DSOHfRLvKiG4rO6
1NGN9UkdG17Xc1aEiCNM2vvkL3kxlRyQKZxntUuPosdogLcQvVgzkKCQExPUA81UdyO18PY+z96s
K1QXslBElzZv7Nhv1VVNL3+cMk9le1CdiuAekPYXMozxC2IcvoKAXxk5bty8F1ubn4tQ7vZMBmSQ
K+YQy9HkWyRU8to/ivKTQeyEkolxy227nsZ+MmNEDd5vfqpxTYYPgI123MFIWeNH2Ngs0RREeCHS
/5UqHwlzaNRYkJXx1MPQc7m8/K3otqfeXRQ+RX4fMQQpp4Nb2qWGd7DS/1iAU46dAOrPHSeYkTIW
9Wb0PJi7xnLMeYHG9jJTq/Lxasyk9Wg4rk2c0/yiQeR6NYVobfkVWKy9gUjORzRCn0d4v16+saJh
jq497It9okxjrfCIIvPerNo/Z3fce2GHOP0tOKc9059hv7mrXslEKcH2balhNb9ODM3FYGlUZ8tV
GjBDJn6hqGMhWeHIU7wQGGJ8BlDgJgGOFgBQGQ9DvD2r/PAyiCR+IabOC3lSR1F3QDkMPn48Z/hO
jbrd+cPIAVXicDwl/xUD6kqUdyUnW+QVAisLJ/hKEZMIa0R+BtZEhrWjDjriEwCpr+1dH6UO4lnO
Skc8hsIfbe5jASVzgSHN3xZXTlUOYbaGvOeIEn6k0Rfg1AFMBHYgk4DUvimD4t5kEp2uH72H7OfP
CYUyIaZ8B7sXp2NSYAtYuFAjs4BG025GWygNnn+fWUchlMMoqc8DDMY+wiMLpy9Mh9wwLhQdGU16
5UgHoBV1R0i7YMGViJ6Zz4x8r/1tbM+G9+S6Y6qUdheT86l4kP+l32fe8Ez22pMbkAWO9mxCMiLP
uGWojrIkK/WwoNgoWU0KkmKTJt+ryGnz2AkrJlb32k5L4lRhzuB3tMWUZEkqVG4lb8W/caNu7WH/
Kmw0Yy9gpntR8X6YP30hhX0xBA5bphmi5TuwJfJcwYl3cZPGQC4fE0UZoEwJGVDrp8W9uZzMd2cT
5NtyxvM6Cs6a0rfroAfN1Hg7HY27DI776BWXiPaPFmq6cBQr2yt+60Wim1ssOoWIIIVn+Ycvzugn
U7e1D7ojHJ3YM4WDWkFXmSptgLCXrRsobrjn2BCVw5PvIGepoAZIb5q4RrUrKJ5Rs7n1DtbtagjN
XcrerKd0+WA2sE1mSwPZxngiSgvDCpv5eY0oHx2Z+60aR/SU5hY2hBhdKKw7ytjxUCUbaLunhY1v
RfFTW1Q7eiWyZRzPNj01VymxgrehD/grAHgfrb8w5QnkEadAnj4h+nwTqocri93sViyGlJHb/m0H
v9Oc3zD6oEROsBXBimuvEryBJJGaS8yNlIW1E9/l/bkLg/I41YreaULNBp/vxjJ5mEqBX8jX1oiX
6V8yY5MCksvLU+WfrCFjMSJEpRn2ppFPr2G2soxUq4yoeH5a9ZHiLrXL1Jx7vfIoSxcoly6a0aFO
TcAlseF5X/ubATxgcHo5lE98GmXqCEXwOrBTo2SCCeDEwGtHF0aZXy2A8tWKVvLrOl4MafMtcQs6
5nYNncnSWkg5rJIqFO1rXp/wO5zGY0HBGQApJuXGfERsOu/bMqbAMVVZ95mmk3GQZ7lowRvuupy8
UbsjltdnbMGCJQw/5Yx50TUn7o05Bu323vfL0vZiDAQFrbtwpiQSwqq0eHZ8Z7wErC8LOoEKmuj6
Sb5lxfJcS/Q1k34gaY0zNAc1QG+gRh/WC8Re5xGluk0ANk3lBP1l64rsQIqrzbGvNDoG0zqHg5Tg
LmK1Z6TVpem9VPUOgSPGdJiuD554BxOuKOsuHh86nFNxDq+7jvuJVFHs8zLTK9uXVhiPOYwCbV+y
jKO1gcGXBBvlFvpQRhiRzXfRgxq/NbU/xOC6i9RGYjA/ezbACO5Cf6+ryfEXTjUVe0UuXFtketNe
jF68T7uV1AUwPVECT9hPR7CzvMN6/93OqX2p1BZeUKcZE0KgKGYF0b5ubJ0U3lzbLi677hPpwbnJ
ShaP0QgxbbSTK/Ak1JZOFuCvdyC2nIpN1RIbwFNVXRQ71TbNzs/eLxxFuB6I97aBvggAPqxPzdSj
9O8ohUXLBFh3aoLHJdjTDoqSn1uE1N+75SYPUcoKlby5IiW/39vZCsHHCHkn6wO8oz0rHPTGLzDt
A5guuIdmRGnamH0uBfINvzgVVv/VGGzGWSdft+3eelgk9BmZNtUEMi/ReIvmaaPvnFYrEtdZHcBv
pFHvZpVXfkvYuYdcdZMUbslTNw0AvwtJrDD9s7WTorGR5xgKmSf68nM+AsZefiZXZDm9rQiL/JKj
x1wYwzEi6rjBvLQC+RCnF8oe5lp1a0RD04sskzsBzuPLxB4LIrt64Ezkp9VwBwwYEkesz0gAIigu
MooHOL1D2vGqL/qcjEE6Ge6JAhxjPDFIxNUwWHToJza3dnAx6IIHDEeIkYCtaMsDWT4wWL3t9rcE
14HINuj+CaGRmxtc2flTnL6XNexB9h+v8Pvw3k/XDChGghHw1C/tw7CW+nSVW5rGxJnmf0+XEtyy
xLdvdwtzLQIUdXmvHUpWlIEtgZeZc9FxBcjwCiHDXxPxfjnQp9OJF4yVMt73aNH9p0XZM7LKRfnm
sKbd4/GF3cylAMfFJiLPxPh3yB0fYSyCQoJjEvnTJX5/lD2OdCCdj+TGvlRXrLLFldiq3pLxzCiq
zJRjVQbqf+GIicvHkcrOmiiVV4FfYhuiA0lYnJ3k8Xz97WdUczct33dw/mOc0cv9dfGk2Qc/rGaO
7AS1E09j9VbGiXGIKv+C0FsjbM8Z+xHcFRGcBwGel35bfIBiYrM7NICNQDi7SAgrF/lxX8sDEuMK
+fZliUc6r7kYm5V0hxkEG3pVEj/CWTTIYAp57z3SP3VvM/ItFsd1lyqEvqQak/v7BmSAZE1sXsY2
efv+Zc+7s5999nia1HoSUCK2k/wM0KLV5Q63+BY4Vt3qB5ICf8FGm/JcPaE214M4GrbjdD6tEPO9
3zW764a1EX1IuWpl18La+goaDvUR5WMTCVOVxn2+wZMlqGP5pCheQtbc4rNPjLTaMKRkXEg59jpv
k0Yh8rNYWT4p/fm8jRGBxFNOS36hJD256SHIP6WWhLNcam0ZvsedB6Rk6BP+YuuMMDDl6kwvPQ6f
4VLq5dnT6WC0KPGoYsYI6u8C97CRMgF7a6J5q8Fuk7kp/vWmGCe2xFU9tcdmHeuk4UNkWh1LOjaA
IO6goc9cLqQITaSwxE2FKWujLJC1CWp0NDtuJB1IfVlcYPVXlVGvD3JGy2v4NhrDU4VN6oL/JztY
N5nx42Pa/HoysRtgw4zrhs6tAdOR2OHIDFGSATt7J2RdcO1x7A1W6cTzO9s1agg1i0IT/2rfWmo9
NzJjt6ILK9JXX/R9l1O82htRXBAbOnNLGp/jG4xDSJmNjAHLYRtvIOesFmxgXhKlsf11YdmcTTIJ
dIDarB/rqWC3UV75u6oZYnsTZAMvdAv0H1eVJxJUCotPYwTgaIi4849pjupu8pPoKo+qUp9iHNuV
j7FDEjbolUFiVP9xurCXDiihr07EIsBxSpojHer8N2U7AeiJRHipZcrDfvPlCKH3hG4Kw+pb/F13
jyYK0bpUE5V+mI4Y/IfbeRjNWAHO9IQ2cj6ZVbGvOk3yF08QdV7j6V5DIoMI6fdhwxpe2/1i3t6k
utWcA4D6uWx3LGknEcUvRK5cmATBNr3SvlV3rAHSjTaVbC+DQBpb7nmUh/jUz0jnOO1cMn85lQN/
D01UdiHiYF7cl5sNc4cVmfvYLo2fxxDlQNV9QznI8ZN0l8nCBou1ftYCBqFafrtLksmvquuKFuee
Lu+FDupHOXoivZcEHXTDU56VT3E6QFz/c3oIi+uZ1jJSpgp/nkmV017hDXQudCCv/VLhBfUEErsg
twxna3EJhi92mjbqm8Ugt6QFoJjzVHBRfI6X4heB4PyhY/nGHeWvlbSgXnLeCxL4aSdtiz/RKcKT
FZHSYFLpgEFWHLjUWLNqM2ZmE7k3XWLD0DpDxYYkokQjJPbvIy1CIS4mzRBYav+VIW5l/1WDF2Hp
eu1Skq8Oso4aaY+flOGlxSsVaJQ9Xh7KRDdPOgC9IkYgZUsEoXopJ0drt7xECfZ8uqlSBuitr8YI
l/7kagZSx1LuRb2H6kaZfSEzwPhbffsKCj+agka+cC6zYp31els4/VpnijzH0NqLz4Cb944R48SI
GNj+uJ4nXBKhvLJyMxQnxcGANuqxts/ckEbq+l8g1qv2CdxFSJt+I2Gih/98tgvV+/xKFsFgVCVL
/VRsdQYZM6/yxODDARP/lG3HY/k37XSlLXrjKtYHRLww5Rexym429ru991lfApYcbBGfLARNNRfp
boBjxn9UVQntUmz+OHrIGgE5DquAxCJqPSUEPlkyt0dg4zUJ/x2E1o506ZIjeeGAMLLDhGA8E8DF
JH5JMNWcGgXwRtLGj5kZfQBqqmXKd1ZRvDctPceuejh5ewmdmInN2/SMP65M7iSeQFIQSCW5rdox
KKSFILBwObfZ88NY+5KZo+3X4KiZsXJvjcfj3bO2KNxLzD8WEZ6xVxQq6mhIBUB182sY/5IWfIRJ
T+mZmdhkL+AAtT7snE82DumEI5D50PuZqZhzvTcWalZ+XNBzS84Fx6AAALIMt35SOEgrdIq25Yhu
e7fZH/yJKUwePeD5QPRrenTFVfZj6tBkasqZnrKuC0CHB6jTXZT9anSVI58fAAhCXdtq64idRv78
HyxdmoLC6d3wwVHfiUnp4pGze7stLa3ggDyLaxworb60qlBB//+QUst9dVsUapzLU95LPOSgXZ3z
oxk47/PdFaJabSRSfedfOZSrnaR+oi2EHUvOwfP8sCfvbwEP62UfZevvp2wpTO2i+PAM+NDPV0Im
3fCwqkCH+r3uWSqMoeR+Gsq6+iUIKz72XNoRVlXornv80ul5NBCdLxXhtbnf3hvZe3Jl29icJQI9
KuquuBicFMJpHn5npjcHHtZ0BAtxjBVoPvdxQ1U0atlcFAvrUUBXuuIYBFek/59mb6kJS4WOkSZd
DxXD3bgTRYjNf+5u+w+zPq9cUQ8oR25uO8uASMHZ4XbH6u1kCMm86FfXTivAf1HuUsidnAo6Vr4v
ignbZ2/RcXovJK/txs23KEPIynANNyTMrVbYsJeOScpPWNmAcaPWoZXZaK0z0wkeoLC2pmBia1Pi
AnSXJMIOi2t/jMiAVHnL06yokqjxoqFkd7PaSCQHzgJ8jS3NjTUuEjXCmep0C4nYO/k/RUIWZzbo
z1l7yaBD35yxbFgAp3rr/GC8rf3hjGgZoTZ5zEwTcMOEs+KwTTgKrI/UutJzJ3NBLVSptr2R7RzR
knTY7hDeKOtnxqSSm/he9heed4WzkiAC/cXhJEzK+plUdkQbtUx17S3EPvcLplTltyGW5sZSTUGx
ScStjJaR/nJbNn7lbDTwLa4seq8AxE3sUs/AwtYS5wML4AAeL+Lk6TcKb9yAtJWvaLHuuFsMZ0yY
zy6/qXqewmPsieYRcbhj/7Eqh2HGmBlzU9jJ4RsLaEL9Fm05GQmoLlkxQBySHzp+CJiWSh8V7UOR
6zvOWDJWio7vZvPSZ+MItnbP18GfohY3EBveBsE7YbPVQp2xJ7YGtcswbaIeObLVAcIyG5ao9d79
fava8+Za+AHOTKnIzkARd/q1V4+s9aPr5kTYzCovGDv6Dv5NQQ7X+OwheAcjXF33o+JSvODQtn1h
lSiZIi0mkPgbNpoMwaR9TrIlug3B+gKc1jUMsRak30F3nPcpLx5zLmIwebuOpKigxoWHFbcbZCyc
IYmBK999mp6EoesFZ604DOJL1urX/iKnfRAI3q/DQPSBgWTJwkbqT3A/MpC473j90Y8enT2EH28R
jKaxQ8fkSzIVHPck6fqQaOlDyXpkvfj2wlo6iW+aQXaeU6N6j3YqnSnNJjNyDZG48Chg+FtYiJCC
06lpxwkkZsyeHMlp1zKcz5OflBC1m1nYvj0h0Twga6mEsE611NXbZffLSbZqtvrDlfHB4j9PfDTm
XRcbjC0Apqq48ETA7axJ68ONgi0D/F1u4Lqc8yKrbui5fDa/XvSGcn5/SH9f30Q9AuZF05ArnbBH
0Pgzh3P5SU46NAyB2cxDZfH0ckF1+MpA0Qz8b5VbD90AYM2G9nbzXNjnzGjtuz0vF4a7No54IfRK
uFSkb3byy/2jrWLVJ9hfe8IOlVjZOcKbWKSV3Rj3EZiY0kPDrlFP7/eilw9lSbzcKoqHDw66MBmd
x7haUDA8qOKpavsxxt3he1T0OhgpyrJcFUwjPjt5RvgdlYajJpsO5m9jwXb16WqUdhX8uWikPwgW
HqxFrQW+A28bpJ39puh0ZqakEL/KEn6RtYspPOdNMabD28ExCJMZ21415IbRGDGH1lsWvrAjeJzk
9jXVnewv01HCM28ih+8w1lnW6u9TFwlEnJVPOiw/4KA+0jvUltAL8vjbeehQG/s7zmt+UiDZddPa
kCeqB5YnULais3u5QgsUqpnMuaeY1N1KT1zlJzbyKg3QS+D4DxWiKayl/69Q3Dg1jXCRewcdnfVc
hkQJKHcifHCc72H5BcCTZ+CBnvSmzHMtgH1+PPZuFqk97St117tC+zpvtTKVvE8A9Mnt86Mt8yi7
1nGG2IXunLydadEoUze6vF28mYaZyasBORqWcnfr2l3yPKkIt9P9EJBBPYoCxDk6ttfSUOvi1WlC
JcZzOvoxRXxMIilyGXLn67wnW6m0d1UmxudiObc0iCt5YssUr1NpFns/I2o65D+naV+SfcV1oBV9
RKSpazGYL8PxmjyFEKeSM+JlWBUOOMegfyAXcZratJGqrLumlc3jghvA7jsyADzIaooTp3aL0PIp
/aDrFy8biIGQ27hDPtWt1ZN4+vu5xkhC/BzeToKZV+Gi7Xd9UVCCZ76pOImbUAnRlJPLGMutr/qH
1b0OuaF6yWmNqsyqq0jZ3JlGo6OMihLOcZZcf8MYX9hmLh4Ad5lowF6cCbxeW+vB8QKcVQV/Vl/B
ItLeE7eF33zMY3nuRxVbcyipWMMZiSV2OUGw4rTdpIF1UOrhqJsKHFwzJZTR4wmStOS7bPqcJxLG
kdaUslP2tM3MwFosh4FXr46SanXiX3iSpxIEZ9mDim7PTqYwnbXJ1J9HUtHV6opWekraGKqLf1PD
m7h9qu+6EA0wjdXbPZH5VIz3dL61FC6nfLQKb14fwrN1FuVicwQhbRHp6D9pcdbESBWolai+kxyJ
RTWrZVHUphA3TboeTRv6ieQ8Gg/yneuQDgXMU5HJLnteUkOiSsYdc/mTELbWELQNsUhWQ0fGLs8l
m7ORKAlRAtJCyHhhVMB1tubxla+hN+yXyhX58nQ5J2JSXQabt0mIGLlu8CHUOXXay+Nm2HHLYxBF
zJUxcnnAXDr6pRgS4o+gH8mZuajkTYsKbppOLF4z90ZEubg6k63CtjodQLmnXazE0KzZEL8Y53+A
J3id47mHeK5VF6JTuF2InYPdAIvEo5Eb3NkSU0VALlF9mtXWp0JbAIB3anMsWMzZODytU+BMS4Gw
5PKK4mFqYSvCtkeY3h3Iazk92KHp9tmLJeDj5nZB9D9ajAvugTMTT7Hjcl3Z3gNh1Cl/h5snj+vw
qw7HP7Bh/vti2c+jlw/QOVTNyYQtjlj4JcRQ7px9dW0BcddqG8o+OS1lRXKczmBR1joajvK/VHoi
sBfO7EHt6gjOCYXMcdfrCmNb3MxZ70zoi5EHHQUV4KhrTml2qS+A+GxPkTTU/fLtZgRm2t9/Pa7d
JSwnw+ExeToAmm5aKOtK63iE6yf2ZUk2d4+VeH+3RvlG3Vbw+uPo5LuovO66PmrK84AUgeyCMh5c
M0PDXH/CNcoJcWTctu0KjImP0/OOaC5VxMi6TzHVWj1iupJOfpmyhZeisIZnsLa2t15jbuqOlVUv
NtjIPDVqfVNHrYH6w3DZxXughiPjVlsUDTgPG0HZlaq8Aqi5qitgXcvIP0UUkSoXLZCW094RwrTF
x7tXqD7GhBDynJmU2R4A93/oz62h633/smAB+zd4rg1GhlFh5vbITwkVNyyoc7iyKbkQSnO0dX4k
ygnK7I4qEa2zfrDAH3kcCqa34JBoFr0A1mwxyrPSs8rKa6MDntCfxJtdCeVuqNK3clR9L7KZwCps
TZbPjB2glbT3m/TmSO1GzoYNs3I7QpVoraoaTZhFO4hl51tVJjDS7/z6QwdmeB4cOmgV6v4Du47D
SbM4BoZ3EM3mbsCZ6gxTDV/pd7SG0TJw2rRI/YFkVv1A0jEhxwID8y3jAjkjFxMm9FXyL1bAlMI5
ALb6muhPWP5T88BHXekhnb4TyO/xLvqz8Qy7tr9YcwL9NsT/1ef8Kcg8+AKWKpZOBiIJypypzKId
qGr17cCGCf4Xk0jBopWNZVxvH0saPfUX/T1kegjwG3tE5ZrAvF0t7WgZJdycseVubpMbf/FhDYMR
DDLCHyjMOO8inz66cVz9XANRspBJlJOkfAi72CHP9oWKehn9v60Uiv0+crj4h2ZrabdShzT/T7mA
dJ0vgd3NxKdl9cyy6G+inPTdCs3Qhc+Xpk2NTFdgaoo5m4pk1rFGxnXKKunKlK+DTtbZySsN7qRK
ANYSEwFDLhS4BaGCdkAN+zYNgXsmv1WNZ4b/OrjC0tli82Z63b+czD3H+xGrwNtEP2omxmitaFTK
zuF2fy9fiqLKB6QpiRwAmgAKdWjMvotNN+X1xsWdb58ZP9rtyzvlIfsgFve5xXSr+x099mCg8ANi
S+gOkkji8HqKo90QiCz4oa2Yk/OVt6OH5MoqEy2DPW8w6IQmTP4j2gzefGUS5JLxI4wZY7XcIGxt
ABgEX/LXBHNkYO4TqPuVhPdFB1vl7ifIxKh3GhP2W3EjkRPydmOAzmPMzPGUImhQT9nOxjPNky4V
tt3ojk6rSav15o3J84rY48YC7TFWbNxwuH5lgjb0MDYdzW12XXJBM1w182X5yfUM5DnBLMKsK4j+
Hh4jdQs4iUY4Ctzwv6PYimI7bTMYuX0gxMkcJYRXr25crV/sQwvgj0exupztmJboxK7Y77+wCos6
mQ8FVRllFhQoqnz4XID1Jd6k8Jog37mdsMfSuUviIWoRgupQf2wB8W6NKzv84CJyrOsVRcsurqGK
ZWcSFHLX2kSv5OYvC4Y2hHgPS9GVO+wL+LAdibAvRJLM4dQNRlblcKsM8ANp0lwNJzWHBY4iS0RF
82z6OAxO2ufHUnOwV1mNDw+B8HXuM8Mwxoykcs5F4ujKHzBNPxNwxJTDVunaGEudbdxhqrQPzpkP
ipMn6VULsqDhRTwqr/7i0A4iwi6TRCFBA9eyNzrX6hxyl5t1eDxWLAZjUz8F1JJIzVoX3XAizktR
HhiXwMQM3m4keuUPu3eRVLESZpHFQ9UYu24H7yogQ2wNPaT5yN/dIM2YxTNeAGLSy0GcYJjWmZti
bEWa/KFjYXiyIXu8ho1VHI9H+paWVB/9Y61TiYRIHOZDEP4gDqITC9oeGRAcbsKrmyMdw//bybg4
4tZP7kPcAJafQ2E6B0ccEtpJY2XFNobRoZjIsjk+Uyty1nD5PX8CTo0XovlPrBl/GdMfhBTBGBR1
eJgzb74myHX9QivF70ox4+Zpjd668rDHWkG6cGBpk3g1nJHBuNFVOAfCOr9IZ5ShnY99wJL12FFh
tZKvpKsS64Lei5Sx9YeYOXwJqTuR7nsMetC9FKpJMT7o4tBPSGpgFFqZo1eTJy9QLCgZ8eKvgV22
K3UZ/0kp31ha2ndqUHfbeeUoW9aMdTrhRna33uo4IaNi/oLxG/UiUTlu1Jy0EYB9ZvmNS+B756O5
nXp7jmNWRMri7zszLF3l9jU+HuN5IHGWZkh7+tyvt1oEzlwUsuNwhfq/2gf58WApVKhZeVY8O29D
hw7i1XtOjSPajEsWatPgq6pe2Q+UHUZOuSL7w3ZZh6+dAdnUJoz9ZJ2B+FFADz489+zQ9QPzWunM
c+xdcL+nEBRt4YETKiJwSLvp71vYvywJ70yNVu4nlSDwI0aDj/KCbAl3FF3ld0yTCPDkXJpNeQ26
IB25BF72cU3C3qnFeONx8rcklBDeiK2wTeSZZFw6XeQkL8YiJ9t3pa1mHyxEWinOvulbiqyzRw4s
j+8jOpYcsWSelM4V1r3uKWKUOuBhkfgFRe046VnTyCzKjJGDc8SnPbk78j06yckwVaq3c3hM0I6f
DkKBa+XNzvvYGW/oRZGZtdDD4VuFx1XSVmEyn/Di2l/Mpn64uiW6QBre1JRZ5QqK8L8XkCpkkJSu
PVCmOqmqIxyRECdbOXBf9ZQCynMdJKSb/+GkHW1+xJKdabr6/nJXf9Sg4TcT5tRC01I+mSrlLKnL
FKqSTrI02mzlByQPDGsT4feIfc0DXBdwU/1CDJogYt5oElbFTcoGEopUDQF4uD3EbTFFbRwF5Mcg
0ym5DOgrvGIH4aiGG0jaUMN0LEIhHad9/Dqys12sw3StrXk41NWKJhcAN8c7CsTu1gG5c+dxfA2h
w46JYB9aDnOCJ6slxOOkCgLKCqdZuM9+QCYLH+mU0c5dTjqo1Iajb+XT7dMurxMngcZ9/w92aOrD
5CHc2nn44ERRkny0ocxtO6+qP1LvyMJ972cBGpLbxpQuLgRg8qKWh2TJKQwXUbABG0xJzY5Wwm/T
UdV2/2S091YXuBpeJ/+j0mY7nNAHlGQRyFwDCxpsbJOZA8V9SSmtmzI9yyhj/f3lO1gUTgFrpz8c
6XH1JfEdZZewa9nbwdFUGG1aSBQiBiTZjCI8z+QKuS6h78iQbP3OEdCLMFM1fSlSTk4rjOMbNAip
+VR4TQbM+xmZXJ7aXxexQzhyLltWZaDb6fg986uBgYI4lPH1T7scvgAXObc14rbA3m7DtMlJBBc3
j4bJfZw8bJCjF0K/ax/8MyA3VbPPKEMoiG0BBOhsAa7juHmC+ev4hQiyc2vEiovmJP2cQSY/3KjQ
+oOtoSKGTJ9pyptoUpDtrFs9ZrPheDeUcLDvRJNiwqMAN5l199bymWfOcN+UkAqAgLPjlWK45Wlt
vkpQX4SXiuUkuWF/DrU1cpgszuQEK+6PfzLK+OnUToENUjT0rZSr0nx5tX/lTgGCWX7HrhOzFe+S
aIL1qGYJSh3BC7ibs/t/5epIivQ+B+cqfMt4cQmDbKLzZhUW+uzHnP4dyM+18SzSl6vW0GTk9URX
jFjMaRaXKH94F4hnppAOjmmjy2pZZ7VCsUGWD6xKwgQmYOIyuKw/beEyzZ8TL1ZSfZYyEDPmnSjk
Zba7FpaFZ0FmArF3b20qmFGoHXnrF+Hhqpgf5wC9WUSnvsg9QgrFzpI401hCIW50juaDhjkXL/ss
hRe3a39sh/AWIk3/JUSP/1JUDh4bPwgDjOZ9xP/BBIlCFXO0aZ0wWw02VO+WV9sx1XpBFNVPMzcd
gvomuQ7PJyNvb3IIPXP6Ym/O7GuTPcUL44cYzpmB1FEjXxnaeNF7V0sXk+yJHybhczQvTarlXQ+j
FVJpOUAB9OkLLxVI6gLgJQUxIJ7CHGOZHEwC7hWI8hwj0TNPISDp9vGm6wvvoRhQwzMEkE60meR6
poSL3gUW28hE5PtYD00GNP3c5fDe9dMAvHJPL40k9ynjbjZkh8ChTY0Brzoj3sW93VLDYUUSa9c4
YBadGj27WKlkXOUugHFXOwOMRbbN3+pSTBQWSpoe9pHV4ugDEsrtWbfM2b1wXJECs0U0WaysWc7b
e+jaeD73E/PHIJKTn06XFGZCp8TR9W6pru+SI3makE3d15hQW3Ir9DZZDuzHtRvIrUvT22tPfaQ0
4D/8kqPSKkbCaNw8SlxizpswICD0ZiA36XW0rnCl+hDjQ31Bej1bSXj3tN3eq55pKOTGF7NQ8DkS
Y9nuzTKJQKlbwWGrlYQZJrk9tle+fjKU1Jo3UeB+w0KEBy35v4VEukyjugHgqSUA8gGgVTFhGPs6
644ZORrvAMIBcNLQY13V8r4VPgKAvvoSUSKnG4kjXtqCELisEZmzq4hJ1LgnkhVDtAf8pkNYAa0Q
dUVNbUwTAAeQ+tu/ST20Fkq3wbN3hAbk+5NMRMkeYiJhhtl2UnNvx1pUFNRQML58orWFSTwY2Yrh
pG+HbEQOvMVPhvIcMTApA/nXtCJ1Mx+yjtc3ruepbbs0r7R4hI0a1CvxEonVEDzC/r5mebsVHltq
TlfLdJ8qW9Pks3bWf6m1fg6Xi9X/rBVU8ONPIojx1TwGY7ADYi60judDoTh3EngE3vqGaHKgdXYf
NTP/8k9VtQNroQE7MbgXZuAVxzSBMUrb1txl+t+rRycwihoFwXrvdT8mE5q5tO1WtL11vu+n0lDV
DfYFhIDIpVsq8IFsDQsr9D9WAkaMAtrH2WuGGQWUlON0V89XN+XtxkB1BRmClEr4Ec66s51l13kX
pF+cPI6SGJkL3+CGHxp+l3qXnN1kxQBLZkI8K6rRW5VkcAcUOeVM0T5S+kFcgW2RNyqdPE4Tu8Ke
ydHkVtrNzWTogZOzvZJfWVKPIe51ua9Bgyt8u3wGbCHmsxsYxTJ+764yxG9vuttnMO8l5XXRSggz
aDSdcUACsE/Bq+BoJntP5iA/nTKLhOhWxht1EYhdugzVOLAp7Tu6Vhx014zkPnMuBoPzSJz5bsPd
axthlANzoDaMnTy5K2s26GCXiS1dyRaQBiFlf6Ivl6s6VdSwUG0QjjmLxoxFVUxFmqPk0jiEHVyC
4JwWwtRXA1XnmiIanv0PF++uiuBgo+pzIidk1W8kHIGdzX0m+ywsrVsca5bObQHurG64OnwA5/jH
LtE77bJ1GDe08NM/+aDdJWOGNyfWebQhFGu+p0YkXi/kU122AB228a7a7Vf4xO3cU02lX79TC94l
35/f3AivzPC/T/ftB5ErDfc46/B2ciJbcZ+AHaxS4QwqXF+LoeSQ0XpxQ+5ZMdIAcwbDT6ySs1az
TkAh0Zco5eq06Mng9iN6PTj4KTngyvkYzdmuoUYY51svG1ZjokHZcRzcYet5/B1Enw9y66V5cfO1
2bJW45chD/gG1ktj8zQqE0tNkbF34kshG8w6BXkD2SKdWAYsqmzHD0O1wPuUtw23zwvkXPF7y3pk
PRkLGb4jYzEi5DaT3FxG/FR2U8o7wmDHcUMBTKqECXESpX2Atwalfs+DqSYCXG9abcHg8JejFE47
awCyvC4RQ6NeX2KO8Y4ehqKLtkO7hBwInPMjS9RHf9kh9admvUWw2++ROcH+FFOLiDK997JqKHrt
ywKDpf/wynJDynq7EaLGKNGa+HQdfRjh/oVaZbCrTI1HrgIQ44lJSRYgYC1Wd+FNCZvdwZL3y6b/
IqoXJRBabANP831oZzUyAnWSLSG/yZLreuBmHWv0Xsa7DSahokahamG82ghn9x6nhK9GM7OPzdYf
G7ZXJsarV+OH+jfKSSgTqdO97l4x2lkCiU0n5IYSU4wdwCx+9LMt/UbtlYI92A/CsjgPAjdEfSxy
l0YcoKBSOYggIqiwKZwFGfpNNz3GoVGnc9FDWSFw384pNS8sx1Z5hjpK8gORoHpCO8kRYYeG3z0L
YI74ABQ4ZYaYlzVZqjGvFUcZ/oZHLSsCGqtoUwKT/uudXjxWmkPSokz+AEmUTZ/IM6QGAYLV/6DH
buqFaAC9bVKe47DC0cB8RZg7JE0l49mc262Q2/CoLsgFQ7YFRcP+uC0jzqhVicJ1bV3bjthxRpiv
VxoZi91issBV/JJAM84T/lkO11HWPr0NDUclptz+H6eBWTQeEENQpMIAdUq+UrnTXlJIbBoWkrsB
b4K3SXndww6D0Gx33z64SGhLpu3/K5vDK91BEJPTk0dn7RvHqxwvKO3CncXvyQtQUc0w/ICQpqv3
RIdmg0j7UAs9OvEp6FAv4fFxIEqDAAWWLZpLqTWlSm2IMWKJIyN+2/wtUJyKZKydkizzmjpJcHaA
n9zb/s9Qaybozn2lAN7pS7pFeqgE6UeJMLnj9vlsJSFdnTIKWW5h1MujNrdwFqGfU1GQ4DBlCRIb
ewPpc1OuaExQ7ZusJPJhlypJLEJYwHmyW7PB5Ukt4qA4la7DBtwmoDTMizWB1iDzi793pcHDJmqO
cY9m9NTc1wo2GsrblhT0utJV0bXK8zbw/lKPkqwJ2rMjrq5raw+u8XMdQqnFPPTifuDYT0cqSQDV
cqJxF5p8opUZ+mjVMGuZY7i8NRJHU6Xv8E4R5G9xr5fGHqG5w3HM22G+r8WGemqYllqY/4egn2Yn
B+F3A2z1knLAHC/ZPoJ9EFKnj28yJvZA7CdAcOIpt02rnpl1PQ/wLBrUa273e2oemu5p70q99qmV
gnFs8IKLJQHCCLsIu0EYLtgxruYmW7QKu8UPvtGBVpPkyGigCdePG7zHP+hNjvmlNuL18uV4+dy5
jwLo9hDMa9U/ngZt2CmHqXJRjarGWHTk9K2w89hf73B+BL75mulb7ry9t3zzmqQ5nxfbQtIqzOIG
yjws76krLrt2MWTftG+aJ0G56oRt+/UWQ03DHyhrknrSCAOzG+xBb/YW6gWJ5Iq99MBX83zHgqkP
AQdKxBEJ7mBIooRQyhp8ETo0G2bmj+b/52ZB0mboS9aKlY8ozfVBH1IHi6ndEnUP5eXAlSROzlyR
zBJmvnXbTW9r1GCGYpWtoVik4D+Pe3oSHTDE5dKmriGFg2s8ruV5faV0+g0V+ZrZl44UhKwmQE+l
MZd8a8VHAGyWNONzAa1SCLnRoJvD34fAaVcTtswLJCwurC5uGpOoXCC7is6DNUk+npSiFTEjSpSe
/b2Fm1LAu835X7rZpwS9Ln57NpPBkdOCGhvS84n7WCX/DShEBHxgsN/NOvIplyCH9g6dNn6vembg
bf0wIq81Tcmz0ZcudKRw1xCGKiTKKTO5a8rK5oIdvA96nsJgTdzy10wvvaAzwsVv90G/Fh8ZJ+PB
+wKBO9hRXzdZtXjTptqG/YWyL+qVV6d4s7GfmxC8a/1JQlGeyxicwhT95Gl5VL0/yfRbmXdlFyWD
MTdU6+tfCjRHLRGW6rXIiD+myT+NTZcyjDo1BDPLXLUoLlbEVeYOAj0//nTKGPsUPYqV9oALa/XG
jO5wUUcxQtbpuMmu3Doin02GiGAeJu97f4B0anF8+go2/jxOjLLdon2r7zJm2elNwSKMKlewU7gu
kkWiSe8KksJOIL2Y9qs8FroX2/7jnFYtgH/aaE7O5BH0nyXDQEoddbfKWkOX0vr1Y8KR81fv4Bee
hvkVT+CflZeXvF3QAVGsPoWnA5mMxpyH7PbN73lF1Jl68tVBhKISyJJ6K59EsQomTKz9OGnKSouB
s0ktpUthegZ2hwrXFojF8m6SOtXpOBe+i3xPL+KgKcZbW5MyQ6EaPKqimKWpr7nXqhSwaOMadnVZ
dFoOPOLCDSZhonqiYfCL0iqRArTg0YBURbZKbVeGqc1oxF+B8RBCZYF89eAEk/bXZ0DI0LIkg+em
ase4Q+BDyHrTQjuifWPJBEDh09RU9yyhdV4195QXrhAr38JPxkhgtQDwD3BeAPUrjMbcNIm5irye
A+EL3NistoVKgXBmJn/hOGwz2Hnl9PdGZseh2bABRrlSBr/l0hTijLhwnfUwlZoYUuN+EGruOi39
1cAbRcNdDpbftVOz1Nwj/n2/SiydZoUPW8/p1+cGuFaWQJT08g29L4E+aggZ4ATxx0i7hZd/coGz
xMNjK7Ai77m48ixwUypfd2aRn3YMFBQQWDujyYVcN1ie4jSv9GHGo/gCIz8sCtf1x+AE2cUPYwm3
vAUFwLVVODY1YMFzmVwajxSMO5uBG4n/UQpoEjxPxaJ0x9mkpvAWJJUUhnvfLDKRgeWZlGTuA6kJ
QVfnC02A8pXUrUsJGz5IWxYCE7tim5hU37FjaI3vQe3PL/jmddKAKkjGexBAFn6LbUcRA5vuTanY
tiE7Zk8Hx34l0xzyntyK4PsixldppZIMDrsC6fC4K2rYh7YlSRyZDlcbQY+PakJFo34H7s1gJC3+
wtI496bn6c0dY19jUPVT5wQNJ9qgNiQ4MHdHbiu+F0x5JBHwQg7NpL+hDWH1pZ/wB03xq4BiAJat
m9RT7L20EdbZGWax7WdMg7rzFIL5Bc4kjk2P+33JtBINsQL65SP5/nnQUWADPuuva3wovL9HQdrI
NV3ZA7PSqifR45gVyrItlM6wC9vjxDGyRQPCMqaPF6wZ1X2lA13AFBQzSLELBTI64e+Yw0rVvFrQ
SCqXW5k0ilO9qDvTo6IyjtMZD5OUN64JD+FAuxTofK6G2HklMBQ0PMo/+jTxOggx1zUmPmpYR7nX
5y9k2oAnzBTESNz/lyzD5UxwhWd3x+lnv7TjE7F27rGLLGl0ZwuKXBv8oUuyAem8T4C5jdlkCael
OD3KJYYKsmG/rp3q9OYEH2coSiTX6EqbW/oIhsqJV1CC5ckJ7wE+HLQt5PrtYlNbrtbe8noGhwTz
PADmFfqA8d+UH1zHTQDJ+B5thDI2M+YJp4zEThFQA5CEuShlqS7zjkr7F7IK1JfB+CWF7wpyIbAz
BAkN2zrEHzTctHHtr5aGKOVV/1E2qbva3bZAdTN6RYnI69HRTrXb0FCBWNkHP/R9OUqiKKlAhPhe
lAAoKlkzYGXWruqeHpZ0biKq29FxTyWpawYnZaYhzUHA1lv9K9dkW0tBYR1nOJ2myTj3bNIzlZ4/
FvLXDxaFpbEu871F0fKGjWt3M673NukBNOQUSdPcgplSP0uwTUEwvbhVWKKzPWwwLQPm3IPbxdcj
QibIIl9qyKykmOyr+n7yDDkh+RHk/EVWu4O760H+BpnfKAJZN8dsLABBKJd1fBkFeuLoRISfIRqV
5z0GRWji6N2o02Pswq7aGU0ZkYrZ4qRCQrjVv/nm+AAH6I9HzNMwHWYwPYM6lboUs0iu01ImkZvM
+FJh93XahOc/wFTo4Luh8oS2rYhCFB9px0cFLMQPhxm0T/S/7qXQE5yt81zt6wWJHjypdOXpKTkP
nU/86zXc49P9+RfQ0yVjZ6tfbFRq6kEFjkTCyJ6R+LQwsG6ja9NbdYnfS5NHd/35YrHlJhnBDjoG
k8pNKK2EWFZTbEpU0CoqZVzVR+2Y2PC5sQSIc6TL6v6e5vxQjG40QRGEk/pwTDpePnBCNhlT/P9B
Hi3jLJFhh+BqCMX+uvR3tJC2rQPEuL2k6/VjYWfye4CLLtZxhnXi39/ik9UX8CcR2hi21zeaLNMR
3b2ujIgc0p7rlbwCAnlWGu49Sqch2Tz/ueDNOJJI4Hz3D9d3VjX8TzEoJ1z9mqzcVEmyiGbaS1Pf
iKD0e2nfkOHw965+h784F/rw3vpxbevQ1rz9kBySzxlS2mNX0jLKyvSp0q14y8HossVFqYgT15MG
5cR+/LAfgZrIRXgIRWSQjsAqGzmXGAzemDeleJacZIIeYUCnpjNkS84fOZxVNBQhrHhMNySuQrPG
c4Y67Nl+2eaawXe1VGbs7Cq2Te6P1SW9Kk9EuQmOhzjWQadC9bLU9PpE21zT6MJWa1F0Sqm4Ig9p
vSguKZgeRKI11/VYFnBnlw3EKEwVxCl0YH/rB303CGexjp1XbCZ0m04faS040B5GuRjjyLBgJhD0
bOk04nDUQjUTrAr0YUK0Px0pIPhomIFC6+GMPNOfEysZBDkjKPBvaX9CevnWfc5FSFcNMLd0vfT/
UcGwFwuVwj+aTDVU7NWux7bVKonTrXfEuiv+/+s5vwC9bW23eyy0cZ2aQWK29sR0+l6riFBz4jL3
ZquPqjVv4tKaJZWDgG+KSLczGKMPHVjyHQ6MeSrlSdIXRZKZRMbS5WBqcAPOtIXpWjPW9adJGaZo
iKRFU39+0aSALdcXa/5DRyJ6EC/TOHS3eDIWk6HiUWgcfLyLDWKJstO9cVfyw7ZE7mPhl+wKXGAq
AR9BM4nqDq084rYWHigFRMsCC8rT+wkrkuTLwM4RRLNWQrFKil7b6V1gaTuFxh7Pj37Jjfqwoh22
iFPQkI+40Yg3BOTjJdKFw6OxA3RFXfaT90FENdd2wNdOQFKMd9gNlTZKL/+Y175VCetFwvOqAzbO
21eWHd817MpPHf8Nb+Icm5RHBwm5k62XhW/1OVS8TZjwersuojIgb1+ZCdc2oShs4eOa07gOpL5H
8iZ2ijwK3vdWnnsT6A/rn9+E6liv9KwA8Duqy1D71cHMhgVnMp7WmLPGjVTt4bu+g51wMh3GDcOq
Et+6mxVX6oPIT493YM7JU7y2DNEG3UsbSaKQs/woiYdVj6rbsJplIy0QpLD8e5JUo7gznw9sRY5y
tZB5qtJvUIWSxElzPEVDDzfwyHTzYBcj1bQP9xeASeY/IfFWqJh7e9bXp4FRYZvmDwprLwT/yaAL
Os70OyXcB5Q1PgFnviEYfqb00vc25X5LS/xe9rgLHYJGPG95KBBTcZwFFZLuIGFeN4LHFCQ6H0vI
ySEDX1vC7DzeF6Jxbbz3aenMojdUMD0YgxYbKh0FvBXIPSowIQNt3AW8bWnuX/lUJ1eAO5RtRs7P
3o7ylYLGwbPN1XSIty9SqTIBXsLFrYK/1zrG3gktPd316IjJVVbSMr/YhmwJece15C35AUGrOQue
kkKku3HzP4O96089WstJHBNCujn2INNilJT2HhyiiRz+cHHrIEBawyH3uyU0rfTUFULkUZcPHZKM
Eh8YeP2SJYu3rj57ILtHoT4MpbV+9yDaVh1khgx1hqPsSYkPryVSCRP+Co8kD+LKFt3y70y/PGWm
h5cIe+yWI0fr8k3Kv2WiYusq6nw3+y8xZm4MT6SKQSvaM8rAOHo9k9XvHV+hoG0u5gkU8VtoSg+5
T0PLj1URKaay+GR7bX5oQd+Ct7EjaFCqCUMLX6Wy5xw5VjfkQK94a5cLqW3tzf5d3kbsKWYsSo9W
TlioxSieCWy8qYjXgDtD0Q0y78PwCY7gYBSrDeM5cAENx8A42z4QWCcY7lUo8Jfjr17Old20VLJP
lvl3G16y17yfszhFLO5kOLE4vebO056MEA5VuGm66WVpgt5mvqJDZDBp4NOcHaMOggD9r2n4UMEq
oNIUsXIpy1Cdcu3hSnCdIf8DJBRkBgj174kSXSQjBP9hcHjkOxEG6ltmX8IzCXp4BDYIim9g758I
TFMGxG3+/HivlLNa4m1aAW3KIz/Th8bWNiU2NfD+OB0pQreFMXlHsIZOR/FNZxVzYFNsb7Zbv1Uc
zH3M2qgqeJ1DETKtlsfIan1BQKYwwadYJHLnGPIiPyg6UoiCH6S/qk7dDIUG+QQFi1BzPV826s0l
jwN8ny7fYYC7c6eAlu0chuD7gsLx9rl+PnPrTOZzZUmiSooM++lmPl3lyeafJb9ebqhglBUp/Y6G
0rchtI+Io52PZpnAcMwuVW65eQC7vrmZaU7d62FaX9deuP7aQG8trdhuhpJFPgY4FwGUR/XdDPQ0
szVUGl7oA4sFmNDRmsb9fHErzVGSDi/P1mEc93epYlDYz1lpw+5+Cpiy3EXJNIzac9W90YxW03j1
tpdNFiXlwsl7J1S3W/ZMFM5kq+h+1RaAgeefWX9nx3Upzmyr8qVjIlHX+y+GS1S37z8HoWLN4MVC
vP7V0pxXAY/DYUgQVKNUP2dXv4XyPyCIcd8hVlH+h9rTD2oRzYGxO+5sN0jMjAfrFOtTvwLaU4Eg
qoQGkBdFYwfVbIVlvrAEyGCFhGwK6SYN9g5SZLhfm0IpCkvXbjwDneURqFzF15hxYNBbeP/AcbwU
Rqx2oHQhHD4tI/C55Uq0otwNj1ReEyGKY/rDNaeKLOfuBjZgrYY33gRW50Ui1U9zfgXk9RParrZY
U+XGU2Rh3XS0M1n7gq8kk8d3Nccd8TyaD7AjaL8wKlnshJj89SEsupkZhM8T/s7bNklInW9SB8oC
Tny9Sv+E4q+lmWEMczU18WJgemzpkoLPyxbvK3zOOpurlrg/AIrMD8phbg034pKrWknRre4TO8pF
/SXjuTniHjiz5e3kTnNCHhnlGbtFeqJ8nMuaAKdJkPVlDehWvCx9bpU2+W+aJPP87Rf2CmhVxBd+
U5UaiY1jDL9mL03mmBxDd6ShA3tTAsJwDD7EOkjxcUpij6f0/eDEbSbRdGasTcaRRn6uKnsMDyIE
48oyY8b/fvugg3gCuZ8nBf8reWjAo7c8tLt7gePUCElx5bL7MJR/+p+GFT1yuIsh8TL31mFQ7/1x
OFa8Lt3tcdJbjYjjWIQsuB+3jhfEQRx7L5Da6qizw6iSIzCt66HmYeWP7zSthz5iZRXQxjhv4yug
VXncKDfaDuQ2K64572Rg2UYFa3Zu0dJrDJswoSJsUB2taGNke1fzKKKqtqIYlRcOZ41kN0/FtGoN
BkgQW3Izsjw6y9blsQf9P+ncGipknLnBRxGRt4TeN69iHhYbKf2IMM4xLCn3HACBZH4u7OILNmi4
Rv52LmyvQq5c6aFE7M1dAHw7nVzmGiywW39KpA7Pz9VgiIKm/yiTzNSGsy5XK5cyp/QAnNUUA9cf
60jiMf/hhMmuigB0/tWhGbmkHNPzdE51E0xZ8T1GGRadGYc2T/gyaUlPL5JMqKc8g9wKpYErHkhr
hl3UDILnjsNJigAsOjyr9oAvcC4jJb9njSOS52aBzZwnHvpc0bBINc0mgMEPomnyq4CkvK6+RLsV
t8lX2o6kKAqOndz7DrSRrAbzYkRRECofggYc8wk/p04m9utHBBgpZL4/6i7YJs1r4O/Pi3YtBSOX
hUM5c+xgrFmnsPCaJujj1YCMxJpZSPRZf2OwZjgM4TmThXfMS3R4nq4W+B5+aJjSh/7sxIUOdviu
Q3mxbyOk0KoFKa9+ezirVSR4IlBZB/cr8NbueWfIeXNDnncdiIEnI/IehgzDIXUbXPAzHAW3Ltn+
+PWmPWkVHySkrCSB8rPzKHInM75UUKsjAkCdWw5xuWa9ziGaVUSQqKqT7C4XfBPzTzAMFQiOhMQ7
f1hOSlroGCR+46ml1npiX8F1ZlrS6w6X/bN9S2zBFXhP2id1cTsY+TqdoXP4VuWHuHeXVO5jNOCK
JOsJWTxQOo/PajDimftr/bpLeDLG7OWxTnTyvrXr6/xjBfqe6TB1A4Wn2sFHcxQ/hBqputqBXb77
dxueBfQDKaFAXTJQcv0hFBRU/vptv+0zft1tI5+2PTKLopFIVVy6QHHy5Z+YbNX+7EwrhEuTTxZs
HFwYK6OIgcG66MSRxLK7ktiUnqk2DBX2p9dqrDE3L6EcxkA76+MxW1BZt4tsNLnQofMO1bOnHBtA
m6UIWJ3STSTQDt2Z0RBasIowxLtseIH7RvS6+RCW9MI/iWbF8mNhMnbdERVBlkC+MOGHqSftXQkC
CG3SZMCwXik3fIhKKGFLIQ6OQ0/2sle+nai0ui5v+jxPzc1pPMtmK6TLQ/KdOTb0X5amMPFsJVtc
xkmG0qA3VokiMjFFdumKS2LENA3wxturQQk5tAJRCfhBSV/hD3D/zexbLXadpIVHZkrjGrAQ/rlK
NwWvB15LPMTQH9ylbXF/0mLN6Z5aneIfQIvtECrpDnsqEwCRKEI8v9MpkWetUFeUK+qVy3MYc/FQ
0nUFfcRo/Zc45m+gyFvokoMgTO6K/YYAoomkfdqCjSV+hRZl/pQIhWQny2LMPAAcn6Kx6f+INXFq
7/C2xQg1XkIeeJD2zWd36ivMs/+8BSD82KZGJqFDMLLNGQ/22l8s3ZoyUY0ZaX3XVpwCCnbHBtEc
Wtdmr9Q1JTJocrq+U9VsssaNU2Ir9ZLhPMJ8/4rEU3fgRP+7MnyOYCMPX+8eInWXaDaYWMpfBILb
fXkb/UUJADtIIsUv6znX15XpScoOGNeq/yh51wJOeicatjTFGansW5ksjlzKhzi2EE0KnTt00wee
PIOr9PY8hjQBLdpNBln/Im5SteOp8IbLcCycSR1FjiLCYF60cbiHCQBvsvwoBC+ShSFJ2+V4pp9p
2JGEQ4J25rFNzJt33cxvEQj50ReQRTw/Rt4WZeKipAUdvER6PLLKdLWL3TNy5Z74DNaJYLbOJI9z
Dou6ykygrTpw6xVvJd5VIu37lF/RtlYMOV2AUdoDTDltZq8kMSN7/5oVMT1EntPmaBmCde/AYmzO
OiGANK+z0JL5tTgqIFTjU63iXKsx4obzXVq/03jE+rxZ7iDePWhT0PT9uKoIRWHTZsBMA8JtTgsm
kg68cekMbUGvw0KkXEW517gvTBIa3wFuq6s8I6SmwdCg2RMhE3NhskKyUzUVQfPexgZ7UpxLXkkk
sEUmlMHdAcJ/Ny7OENgsYOUco1MZAicpeWjT5i7Y5t7CXESikwMrzE3+++DHXp/rkvSWCz2haha8
2g+/l9Cqa3S6hWTVMQ49NJqrB4C7irlGrMI1kk7W51MQ0JIcMwf/SHyGMuQGCqLd114DovAAIBsZ
giZc5XqtA+GRipVY/lU8ckEA3CTUHO4coNszBHvVzQkoxmb79gpKW3A3UzpEzNUblQb7IYeYqluT
Eah8kBFLiBD2VJ+u+Dv6OoYGqW9OmTu5+rlHMkIKwCnBkT2SceK1NTaQnzrfvwy+HF3sk71outCM
OTSCaCVNsgLlt/yMZ/yBkaG9Wo/3DlSfWne5wC9HFO29h6JS8YERMXC1d49ayS35+usOAiFz9pKa
8A9Iq7CrdcsQoXumfy1dwSo/sPn3IaPuiaQhnJb6BM7v7X+LrDm2lTSSKz5S7Fos4rJEIwKC3/Vw
fFbiGxUWswm/E77QwSRiI1m6nXmeEHEBl95458hfcPzRQeTt0KCl6yM0FdNoBrrqJYu8jVWek2yD
qzSZH6OHpYuK5I8GclJa1Y+fiNxlghRw041HuI5vXp4RC7tKI5oR0vm8zRJ2MxJHNoI+9rovIS2L
u9Fd3Mqz/xFWSj4KGDorLGr+iR0ajBSJyyYE/JoIo3ZqMJ4wDh1g7RRTm0Y5jBDZza8J3VEiiAz5
4ToAl46u5zQPZs182Wy70UKCLoWFui8qn6XfsUzleSfBbXfLG5jG/skW1zoCNc6aaq4QDcuyhRjL
BlB8woqYhGOjSY0goZTkYPlzDkqt72Zvzqp8zuoqPyLiUjwhSjV54KEx+98TABNVL5XUwrquWVC7
CHIwctFSGVZYsXjBAGwxwnSGAgIL6etGXncLjNArz/nyOMIRzHQ4F2rNfy8fKmt1YTeDqWCnx6Ej
Ba0wbzq6GPEMvbeXLWmK0G+0krN2mtCs0/kGHk603hvcvNiS8I2hrZMiWZdlQhS7qH7wWwedWGem
dieKAnjgIyBrwWjKGPsDwLPo+TPn/BJk4LTGcI1UTqhiV4NATdydFoS/3n+LCToyrtHZj6iwom0n
TzJAyLZYeBLHOQD9CmNB6ghR/fQsSPiHcsVpOX59K9CZl2s79BOXOLg4W7oTp1+HpjTZ31yixgBV
bUFiBYDojn5QFto6wc3EnO9Yu6TuGhwf8+RswrNGGVYajl35MG33HGbmb3FRIB1HHKJ7tYi6JHzY
2sS+2yj02Iq6EOlrSZczR7ssGbfKY/ux/D91TIf5jR4grY/+GUiR946zB+fOguFe+t2Are1k8Ixs
9VrxRoWDozcuM9n3iI4+N3z6zumP+566+HT/QTnpuUfGJ1BoKJqWMaBIhiZ97Dbmy7dIHNU+Bqqk
nuIDz/QZikeC7pnHQ7wDm5PRgbBVEWJWxYH1maNhcdsFyaVDgGmZw6n1PVyPcE8OuhO/FL1XBzAb
u4eOrJnNx4hashIWVGZqAhFUN/El0Xp3Jh6POS1dMQ0SRsZTsxBVFT2QQvadRqimAle/k/fNWH7w
YvxCnb48zakhXROuriwwFGgy73/ap4M0/M4EAKKFItqjbjtCqFvqWBGA3EMSCfuTFTSWwHEhBrvw
tsKr0/wY+hC8ApGxoq0Fbe07cWvTwgZ9yOdN9mQoqC4u/fdGXlOwPIE43drQvPEVAJgM3dBUW7FH
MO0pqNlrGpgOqpdi9R66gzTWdATJmJdJcKUnUXeXDNT7I2iKSNbv/qzplldZaCgWo+P2Q9xe2ESW
JMN+t1peeboVYESBl+hf6ScO3eo9ir8r5Xa/nnGw9E1vexns3ZMVY35LB2Q0+kmIxrIyshZtbPIP
wwE90Y1Qcm4iDK7QQEORdB0qqWQYASp7Dnd7Qr6MsVfRTJ66SNmgFSckmmPFE6Jln2rb/LAU4CrO
9lae8KsfOr3go3ZUmyff/00UuZtLnOqxSxextEuSxR7l68+J8SZMlGN/7wL+3JgdqfxyEZZ+CohI
JFl92skrSEzW9Ih3WHDtwTPP+6XksbMlkxhFLJGJmYW+rRL6FgfWvTU3H63Glztbi4LXbC6rk8kd
aOT/r/jIgCA1Ei5o/8/tAA7tSyR+Ofke9ruftWIvDxNcmG3NXMCF58PakHyhU2fYS6MjRI/QhQz4
31625WT16MWz2GOOzbGiRM63bpxlsiQCmbkEr2uYudeRoHLISC/eb9OPnAWlBxV4+F2ZwLb9UtEd
N9rEw/lehHhRccgzfVJWBvpg/Y8KsvFjCSHCg3KGXsrw15C4LwV9VVq28qNRy43NIA+nFEXBWt3m
ssmNsSM6HG4JRO2lad1k2g8FKOVvRztMid9BXCSVpsI0/d87D7ldWCJDmRlIPUS5HSgaX71t27KT
wXV8oebBtqsQE43CqMamGNXhpp2XS0iAE0RZrxm0g2dPu06EWq6wrcxPY7dgBP4c+j9iI2kVUImt
AcpzdFfpK73HnvQt6gpHX8t4GYL/fB8PkLI4qE8ECja6wvNK8P8LwacOgLs1MgCD9CfuqrrPYcxX
JcJN7ZtX/qdqZHbbNo5uQMb09lkkVwgAdqkhnaRG0FA0OwqoHWnFnTwRlGzhr14b1l8CJUSCSOTU
HYYdsG/frlbNdF+16b8PWxgrqon/mPyMqSGSGfIBOD0a43xSASNTd+oHzAIbCTg59lm6pYIP/vHn
H9MWr4t6p1XJ7SGF0cjE129ILdF0njGwutFpOJlQfoV7o1EGnwQbyhgV/NledzQNm5pI+yPg/WcA
x7Vqs4ZiKxn3L1o23ho65lLA4YdG/OATyqTpYSmC9jaknEt3LPRt1OoJgJqzxNcATqKSTZ3SVBmX
5Y1L5y34bVww55YJkHb/rq/js8o8l7zM5qLcIrCYAHpdtHeOiAWLt+bAeZxW9Ls6cJNRYz8m/lKq
89FJ2+lmSBCJkj8SdHzJNBHpeKVcOnpa97Nd2DvQadM2LoTYJE0LTz/TPqKaX+oYoVcvM4m3uTBq
3adzLjnx0R5g0yjeP8kRQZN++w25P1+SNzp1r7Dfw+hXVZgPB5f3xmUGks0us29kmIjCM1GFp1Vi
l6EbRVT4PxEzk0f1FdHGeJlzF0x4H0+HTEy/ets/u6kVV/hjqQQbqTOM5HLXyfLQ+vqJQzSvRpl9
L9rLr5Kb++gfsCgfI/dyd8adR3NKjsZH0uqbzMKNz0wuS8YqoqPO96U7cyYGiLV6JEUEvY94WJUj
3NYLDCGkeAfIOuUK2CuLOhFXz2UOUIENYzQ+AfBM0Rs3AEHZmMl9SAna2wWx/GFOaYfDLT4DiG27
qp4HSUOBABVCKVdi+syrnM+YVJCMeqSlWiv229z2Dm8Nby9s8pxrKmN83Rn790clRGUBBPCmvVNs
5lNisKc24X4c7U0UsUQ0iRIy4zfR0yEXPK4QLFXf99TSW+3VW2PgpB0efdJlCvt9DbOH2q8mm/1J
ZsJ8K/2OSvvcKihy3zp7FPof+J+GT3ihIbBt3nFi2vuhwGXHBzt+X0c6+TWnZG3ZnLgSst9ottLP
eewIRkSMK5RshyEJmJ+rYZ5FiCezsU90K5e/4r95B+oC9mEG5Uf/g2Cs4/G7fZJFyZn2JAt7iN34
USJdXKy+GobVk/8lXmZMSy145Lj8BRAxB6uBQHx29geRxNWXSSIl4ygILKbU7G7FBvncBeQQz7ud
gQ9z9aRN3Ei33GTmWTuFrZ3UbnTAqGADcxh9lHS89yihIyHBG7rxWcja6exWG8pgl9nH8MwAl40A
eJEqVfqtntlqFOLGt0F2PvN15t/CaswHRttGyLiT7Q6npYdSiX1tM8+bU7qKRGSxP+FuOXJbPA4L
8N1hSfm/5nW7bow5FjsxzZ0qZtLS9DMaQOZQVv9dq3wghRRQaRYIXGmLqjQA/1oH5/Qg9LLxvHpU
sns/Sxbs/R4vkOBFwxXJvhMPk4wBB4KLLy57WSUifSKe4WZjBN+x8RFFk//VZ7fmYgynLBcpXi0u
LMpPEmRMQ14QcG0G0vCWwa6atPsIjF1P0eaBHW7rxKWmUwd7MrFaUDae4UEsxV5EipNdb8hfKo50
/GzHV9QnLS9im791kP5Mlv+6sZP3W9raZXmi5kDMs8DRdIdpVnVgfRbfwStv8YA3lG0OSTXfP+VW
vomXnr6jC1bTrHeCU5fteIgP45cB+kwqxKVKwEN2SWEfIpyYlJ/ZoQe3CqKstIAPFK4L6kN+LTVg
TIaJ5v1IqQQ1RMoJlzFm2ZvnZDuScIb0H4K+qX2DF2ax9/4z1V5OAUOj5rAc1mZXlPC0UxMWJc8C
0SH1GfhfcGewp/N/TQ4a2la7yTs+G7bJcM/3OUP04TZc0vq7a+wN9rWOAdR6NopwTW7y3xN56eG1
vOd3R83BOT/zvfjDNXCm1ad19r9KciVmeDRK6oRrIjVD/J4TnlWXFWHKX9uRSWUrclqhruVQ5LR1
H0R05nv8okfWry9V080mcvEQ7CFllTDAJoQv3HESXqkhIAHiCtHmGNlMnBrXN4Ebm1jdBEqxVA/z
1nIUoVFKHV4YCJQM9bXotxTJvJHf4RhbmTi/sHSla5QiWmfFZwp2x0yBfTdGXdmLuhGhTI9pTSEB
ZxhMqQ1cYRblG3dw4nFZ2qXTpn2fiV9Li1vgHKBkN5aAJgp++c0sWe/MoibZudGVAqqyc56Bu4su
u5yUgdC5EKUY+oRVsl6xlYNjo8NycdmuGfkHnWq7TK9zA3dx23t8EgvnAZLXbnwMwWfRSG1mgg3h
bU71COc4uQ/TW9BL1AFEOLQscOEM3rPkUzuBEDuvVlut4RIE9mxB6ZYNkOEWgvh1caqa9P/+7ZHr
2CV5NorU6ew474gfk+friqnl94589yVrXRqdqB0OFDYI83Ri3+uScQCCpwqfLziUW2irhPlmq5Wb
UUdTtLy7rPjB8xD7BRi4pSETmXPg/L26buOsm+1Gm4WsNwQ3txw3W/dfZKWQtvH7oUmlI5JbUIac
XCmxcwbHqgy4yk3ssHTqa5whKNJvgQCP//lmK+inofD/C93FyCK6smC7jn3voHhXd+9BlQITPJWH
h3faVBKbV7QDveVpzI6IvkfEzzE1gyicypeVxuuqbHuSLhxb5EJlW+N1jvU1g3FRif3fwFTWu3HN
SmOo06WvHKHpL83iccp79g/Gt3IYcquzDYNACq71pYMBP4pLXkEbA6aWzFinaHFrdrZS4CC/LBcu
mqvyBC196b5tOC2Snk5nBonMiOQEFejaQPTFecVHD11Aq3gyujKWcc5duDXjpeu3Ju+Me/WL+EDa
On88NDc5QXFTRZBwZpXTMk4JcReNG83LAf7AL+KZb/w87FkNE4FK4BwPMtQRS0NRambj7h1vbRlD
rHMdjt5Q7fsWgj7f1cG4qnSG5zE8AfqxtaFulP0cxVOGI7pEm8GNxfwQI8T09Y2VyVNmpVJIvMrQ
HWJEmppw1Tp014a8uIyFbIr8TiH2wux/LbWNtyOOUyXt1VROu+MHL4nRRXdGgvIS7r0YpTNJCf21
4PhNCC7habzSoPFZq1pF9tr/YjYJh8Ssn9urPhx3c2TSpp/TdHjDQbW4jbRBI/XD3ckWLtmZ25dB
gnVQf2sUf3HQXOk3zRU7GsPMb4d5uEplxj6tg1wqUQ9buWMsv5onfgQm6Zslm7Ti4R/ILXLM4L+n
nyO2CyjDuroh4CyGxEEEsk/BjP4eOLZxS4iUL6e8pvRvwiz0HGaZ5Sm+DRZ4UgKd1DvJFXJQUe1W
ggT4bRD189Y0SntD7vzdXpCWnfTph/Km3C/jCzr7CR28WObGw8QzrIohgcLCIjHRBS3e4hTpzTjn
8kh61CSuWa680bLES/001878q0cCdoZLtCYfqgF+bflvRbDPDJh28H5rZMPqB0oF7zQ6TKZiJlw/
FoZBZjEoly+DAzCQW9Nj52UO0g/Ql66xBYH+9sC+eaMIHhFE3wUzSEvSv275Zucg4uqXw7wTgwCo
dkAdVbjszChnrSJ+Nf/LocCpO/euoXQCVGC0w874wtwEjwEySZLSHhCmnD0kBupSIbsHPo+aGT5g
e1aXwDfvKcPu2J17AceG65Fi/A4PAV14LOsw7RhhxfAjoeoHcyVuzg5haLv2vYNAIXGtZFqHxjqh
zsyfTYB1TnrNqbSjVBimkpTFxtWu9fHdtXga1w9qFccDMancswyDG+jF/KTzM1aD/fxusPhgb+Kf
+hcm9fZNPtYd5bZ2meUFHX+c+2nTTRrbksd08jKf4MrFAb/0a+EY5EfIR8VpLy863FJNqIBQWlvR
yh7L5Z4FsRnayioxJ1hDNshTMYYqAPOxJ5c4AD9w7PvX8N46Y7T9xCVzz5mkVzrzm6eLFJvfKx0/
AMXVFtBl4cGXXWIojy1Ce5pylxn3IUH7hrGtr/4HrVY7N7Gm92DlwmJS3AqX+j9cui2pRj0BxavQ
XIdH1RzCuIT+qZRqIWuoVvKAkeeg+Q7V/YlffGVtZdoUC1ER1GcGkc9m8UhmkyqxsuQe89KvOELQ
okU9UwMoeQVOuV7zlBX4/u8IRBxO830vfjILzaC0B8GeCdFUamfEERh8qszVJh4ZOiVagpxZBnU/
IPX+yEbqt/RHWwXf0HZnsDDm5hRC8rkoe/OMmBELsqt9mgN71l0tkifJjbV1zvGfSuy2ka/mDfK8
f0PQHeYV7qEWKOErmTOlxy27Pkt3+jgTOt3Jny+0gaFg1RaNyOkgGGqsO5uhcRVot4hi6NTu8oAG
RlXCfWkHga91P4qPH+taN2MqIjxlABZQPEKIhpzslx3+ggRJkEx4n4lKNoqwYng8EVyk6ovZ1q+e
50maaWCtT47VRR76oUowGgVF5og+PiplZOZGaP9EtV8OScGopRYyUeVUcTVJyBtln/3ZWIKksVMx
q3sVcyMijbOZsgvxOMqQHP0j+zubdeksXBdSzl5q5r47MSCG2Cw3i+iTTtADBIkDTQ0RslzkCv2b
1OvBFEc9s+W3mYK0JaLkM/ttaPYFSnUcM4aJMMlDOkxEh7qlQy42V7XPyKFD7PFbEXNiv8Fh3bEI
6RfN0h9BsqiGfVLNIiVHozXaZdaVg0cKNkEKgAOf4/Oqp8Rt7CKgkv50GhBDYwuEBp8FvGunzD1G
BD7QZR3Io/pUL9RDC9jCCj8TCpQehTwHkDrLxtL1Yauet9VVp6u7DO1kTod/orPM8ozHACDyEJh8
9uM6N8402e704XlENjOOwztXj+KpRkTorMSVwMw/34SChIvfsTLDF9EZBAq4ueeZxf/yrtXrBXoo
IKj8Wz31WVh7BKBFBEjiqzLUI8sJ5hYiSIUGnUhuv4SZJcX8Al+6sdFqg5GZ4SjcNONpied4AQCG
JMq1RP50KxnYkJPJVExvPxTb7mN0Oz4ghu0UBL9BxHm3cn6ihiZBMswWSBjsDWNah5WFe6YgzGjw
myAgCGZJK/OvzgO/arssL7xzGsrM8vtIMVvlF4sdfr4IqBhYmjYSgM/yyd7ndJjE7R4Qs7jA6fOS
5VO0NGibmgkUVKbC/r7XpZioOGh8aHRqIPbs2ZpgRtkViLjkPNjKFduY7hTxaB4guAFQkaMkPxIi
DznRLWXSBDoQOkraNPp6dCcH1ptCDpR1KpWl1Zq/SLR4mF1le5RnwX0bKweiaRu+r52Jkoi0rOpK
tLtwcC0Kf3vLG4jGEIPjB0UaYLXIRimHsR6BgtwRO/tqdHU4I1yQqV+N9jkWruC0jpyZX4MAYoTk
fBIsUv0dWvw9udY8X1/Xco8zh4slp9dIGpuAwV//JgTc4EHbB6z6AGZOyTStHlp+0DoFQYutBY5a
e/seQV8NYoVnisrxJ5k/mJYbbFOg5MYNVpz0Hp4YDHuQA+5bMvEY8VAmTo15OeWw64BC8YMHN895
+3qBV2MEzJqUzb7z0hgCYU7PZJ/AimXxki9hr9hbYKoOHHavL9K/oH5J5prL2TEvh6gz1MNzJZeZ
C26E6C+U75ZEo3HuEbEIHhT1uWyyDoj1dK8IVZ/GPZpVi9yUrKJqdUeHeSxhyPSlhDLs9puPRhor
L2HnPMY8HZK9mLwrF6QtQt9ehU4Few2TodDppeO4DxSd4zI8eD0DcmvHNohnYVvG+rWH2oJm37Z5
5XShhiOigiQOtV2Y0R0QMTs8lumTg+ZPFUazSrUq/fC0kvi8bNwkZ9KfgUzmc/2nCxf2yhJIWFQo
V//y1ehQmrQFpTd/bEOma2tL9F1iiHMnTSgarwA9F2dhY/tu/s5GQAromaXV3vAM8T/w8E0dcnUN
4JOgo+eiGr7Tv56UK0eV1SiBBjKX2p++kAWITrhINDauBOmRbZNjWpwHEAkXEsPRZoc0BIW51lc+
RKbR0Osa61iiP6MJgVjb1QIcO9gld3bXhzcUHfnwyssDdpQChpRhCGkhBLBRbVQ7fH1GF2qJHVLZ
ZHyxEGMsZVvsw9nIo23WLTuruF3AselXAwkiDWfz3pWwAnLS2ZutUFuyrZxTXouodYSu0QF8nsv8
Gz43hEOBjWOBuTit0cM7yEpLGe5YhgKuRxbfTf/sGPQT5cj5JD8wNCbB3xwwIcyK1QloGsD7Jbpy
UQLz4bq+u3oZclL1Th6D7zc4txlKNkwzJEzu5C2IUOiWyQ/CBSPcOVUzi80uTLekzz5GS5G9l8fG
N9Fj2EPeqKh1ej3qkK8rjKcoPaXT+rIj8FiPOCyrM55EDG4IOBQPNukE6Qx+vSTOwP/Ln+7gvN4R
A2Doe0QEsiTSX+S+J/LoA5SfuWCpe1LasDTnrQ08A9ree5ebeTkhfh72c5ibeBTTxy5b97yuXsUs
9HljVbLCSBPSCz7Hh6/WSLiJzXx8zLgTfNWW1IxN0bZDSl8/IRbg0KoAF5HjexyQZtU205eDBIkB
itppShuZgqy8LBYJbe88f/amzpqts0Nk16w8UmoC0a2zHwbWOeqCLQu2657nzP6j4K3zZHFUagVF
VUstAYjyl+mo74NZsti4e/ZJKByBwLe+Hx49aDyot5jjbKKOHOfFCQ9JgTIuDZgW6TP1TpV9VEvj
dy11Shsr0qC+QWATo6UqXxiCGvsLpFV455HsAhZkkpCpIzbPxvDSbqkRNLsMYRzYYKN60AyhxiE5
Q8jqDEqUMsAuINWvuSueoJ27pdjj57/K/zsgV6Fry7B7q8i9ov2E9eOf1lAGKT3eUUNWhk6Y3Jp4
FdkpBq+VmInZ7lMPa6WVOQPhmraRkgXZbHhwH9YVDX7yHZx8MoQCsynf3FDT92qUF76EUzEqAOhi
mW1fnD0zNklFiaCQv9Y6t9jaiMDJHPjK2giXPadO+if3psd1PCTX9pJ0AtikL1wgluK0tT+ZL5Wp
Lpcu2CjjB1ogSbfdm+9XoO9LNGXRG1IkNnEKTQk2/c6VW7uJbC9UDi1xU/U16MEcKjSvAmaQjfIT
VsIWBcSSLCA1oustjZo/MWsFUYL2S79IZowasYGOxZW6Peg+Uitk+LXnwvJ4I9wt5wBsMiuO5+VI
ETI5ByPW6xMpVkZ9hcpow8t30HuYre8w+VGwnvNo0ztaoSm42CMShVYD8U0tKzBCq3Vm5nnlnRAC
b83UzLKcdHiW0ZbAyu97hHsafUtFpWdvwgTEeV+Nml74PE+zuCHMAgoWUw/gzGoYFlixar1B8vre
b3/KH9BkPb1pgazymvFkMOkidt0+4qPgnQnbJ/j9YtNq0lhnVhjvqkwFVz75d3lZ9Q5N30KUWWFc
ZCfzo/ehTtZjdvP65z1gWZyzuV11p/N2748o1iox9bGp/q47v8mQvceh6CHMTPssOzVVhz5BMkcF
AHBPwudb7BLDvikTPrblcsUmvRaX5wlc7xL/tK7xJY5vPDlhtiLB70JckQ/WzcJijoRniDefXeeE
i5KbTQGSno5SY7VqPJNgND2D/UCWINGZxtTMQEwmwKrIfO/hSAuP10DfDGBnm3gRnJGSfFq5rZUW
k2K9cr6M2kOGsyTFC1HQN8tyoIY8ECPNte8hP5oaKfdVJ7XA80nqby1yit8Hw1MGg0AmNhk8t18y
NNLNiGsdGMhYWdfxVnsokEsT1+OOYRkrUire0fB6ungWz03cDD5iGOhPIHiVa25qgw/ZoQiXEJz3
LqkMiOVxG1S4SMKil99zCf0DKqq0xKCZPD1BGPjjQuEOahImPYmUfrTOrQTAchhNhpfhHVrCgL/+
6TzQkDitxjxbKxstw2Z9iC/KkSNIC5uX23yvVRne/ZzB5w62Y/4x4qjJX5yJ9Fgi8/60AhXz4qzx
oje/WSm5FIxvzDXDKDD8X8z3YTkzgtegYlef0l+4UzigQ2ve81W20TS4uweFR37/faXX1rslBUaf
lZ2ad948Y72Zq0H7hU6n6L0w25sGEf4K4JG5nWoTX9ZB0ooSTx6lHFmtf5upLztA0WJ8YMvfwZ8u
pO7guzfMxUaGZ2oAUoElJdQGZiDb76WG0QOvDBREqOqoBMPX0j/xyAB5PDHf+CbOjcmdj543JQ1s
H0bVyNVrdJdF+BUd2sGtSg+7ibrP3BPdVwD10vnt71D0tjVkiVFnAqk63F8bsVzyKmaPt+NxhyP4
p2hJTIhAFRRTvhzGtmxJvRjnwpSgA7bGk/zz3Ziy8xOxf9cDtUFfhsmXGpmZ04AnN1w1mxqt80aN
G5iYRnqSHH1cCprelU5VyaLanQijX3tXX8bOscDCGrvKPVhjpLc4nls37HdsqvgN0xe4n/KtmXip
ga9mhflNzSBQik/Kt9cBhq3w9lkWPyFn2b9HYrwaTPOYdPKmPQoEdIrA3ogY8L9D8QQfHla62c7B
7CGaprA+h4YwsyG9ITfFG/PYq5fxwKcnyPDE0bxOaxU4ecR5HaQUOAPYE2TJDyvnEKfZY+tJDX5i
/3aXXIZEJ1+fS/xx8z/YBhlxQpDk18qPNxgX57xFcJ90S0leRgBV8CHLNR2ZTlgO8eh4yzLFxTsN
g7aie+PdTpYa4sJptzHNg+ABxXfFGNA/K2FjwyDqKFkYfurSBfjdFV7dEbSpCDwXCb05S5O6oEHP
0rqgvawsZVvpbsenOPVvHc7kBeThp3am1aOSbTBslvSmYG86d1lfG8bI58aeqsSJAqGL7EzBSkmW
1twzg8kviPTsB78hWaLTddn1inTFcVIjaHnJmzr6XTOOaerHsjZN7IW3LDLxYLRDkZPxv7Dhw/qs
HvakME7u26R9fq4uMyqxa2yCN7gbLq+LTzNnlaIxczUg4zXb2oIYCalz45qwbiI2PD3ln++L+Tui
EDcopVluSE8ipMA7tUvnyhNQ2wzhaMufSDvS/vft5h/clKbuY3bjr53TIRelRXXvjwka09KUV3vk
zFQ0VN9YdSLoOpyjgkXfKGA6YOMPYHnhbqsuK8d/CMvTLVZMm3Zfa+6/cuR3fTlhzpCQr18iTKTQ
7CNKmgg2orNqonJBTtEvmKbRhx+bNuakoAnTwE9kzG6Fg+3oBnnhHkhwUZKSqbT9vNwzWbXK/13U
xxCp5DnL/ppf0lGh1Ix6mldt7b3GebNHoRYAK16+3/phRYZciZscla2eQ0IR2fryiZ3eHXvHUD7E
PVuTMpZ7W5ds9A2imiBZkFGp4uyAOEWuahxgXrQ0v05KwV3pAeT+kkprKtb5rwwia/StzJz6UBk0
tFJMIP1GwUNsO1goVfm2yAxKNJKLpPj3lqNUaXEKX/bFlVtvivm/1XxKQzlpJFN1X1OEbiFP1DVt
cYzo4h+SkjfkhnMaYuCCnMKCwX4PQaaT7o5PzJcB2gJ1cf57cuhzEYUFbD+pgiVUcVLDjG7G/o4F
iMM40ltJVYvUN5XM6esnPi7hv57VBJkPdG0MosGeIczHg4IgF6n48iwBi5GkYIdcQ3XlhA/amzqu
E+RB6fDlwtYzO9/y49zQIZ83JXHfCnkb3usN7q6T3rh8n3/5I50oAd1OHcYnfKds4jIutQytjXJm
5Fq1GVQeLDwyN2/OLDvERygXBH7Q6vnJEhkeNCjWJxovosPJd0UYmwLq0kgsCSAuAOgO9xLpjiCR
FLD7/94ioQ3CIkaaveGcs2s2R+bVa94mr1vX/OZD3PCQ33t4lGEdIlCGPmRg/QtJMrMu/2Tlehpo
Kt2NIYg8DuTzJZISP3sSwWHQWvuw2SlUk/YwEDb5WT4Pmd9ZGQjoJ2IvdJtHHamFRvpyC1S39j2c
VEl+VSeKc9T8LwYNht3Xr2CL1DL4/8VpwH9nk4vEv94fCeRTbTTlF2ABImKzsds0W+NRR3Gtw1ks
rvWHOaBsMFYBcZZ32sreFxl+eqDcwxqGOpCk7LOtrxGtvjV6XNPtDOp3k5rd7qxCcA3les8kJYr5
Q2wEZ2NM5O4kuqzSpwt6izA2TKLjudDgWAo3c/p+eqxvSjY9JZ49vXMFX9L66Ucs5t5hud5Zu/Bs
sRGIbnCI2RySheLhGc06ax2JYtABRj9pLQCPdz2dR3jW/Znx6lm5Lyfn60MXU5WTX6qNvY5LgpMu
fdF8Dn+K+SQBXkPURAT4T3Cjohl9Wm0n9vk/K5BjU+pbPdNHHuvBtRjHvAV6bQbakmeHvmgoYGce
e1qwCI7brthT/zTyXQzpk6UPHYGE1tDSDM83Y/8OaeYyDv5yJAdxF0Q8fybRkIq8fMnxmKGQDfoW
9I1Lz3tj3xi2D3FDQsZeYImJCZPLFZvvlo9wJclJXIW9kWpAExNBy+TVihS+QhVpwF69rg30COGt
RAhs1ykC3HQ4Ju3VJSwbThJp1KiSOUkn6LGtlLsXD3cfOGkmUghCZkuyN1UwALfdSzKbi3J5MERv
HCWKgGOAm8xhiIYThR15INno4f4pbfRX+SIFAt11rYRW93P5LV0K0RRO0SrWNain7ri5JUeITNy6
+/m6MlCZRNhe7yxNFRBozw+tE76czyDQL2pUVEVLMC1UUpPbjYdxVYWrh8Im6BgGnMzL2L68i7Ez
SmeNO+7Qp+YqClCnxo1bo85orp76alPB+tH0ErDjBl0i/vXLsPvpe8Ph3KZ6/RwVWSEy6FE+31aj
e+hqeapuatRAWKmv+6ukU653bfjlP5HfT0iFHzQyUD+1KR/X89m2+828n5tzinzfZ+ofyrkFAnQu
PgHhKaZzeh4bYkUnGezMWP9p5PJt692I2QF6dP54bkw0Zivi4bnPbQWeiHMZkk3vW/3Ykk25PH6l
OyWj+sbQrCp6SltJWrmBwLqeNYdEZO1hQijd9qtyOrWCptfVkEYr9lx6mIjlYowWepEZOsnbwS1s
ef5czMaOYMj74GKIihblKWUtjJUKvLD9Wa6Xa/kYNrDHWOes6fOHeQNEUcN+MDdK2h18Xqncdy65
4IXy/WoKvoih0/hwEAmdAp3dO0nNS1cXqOPZRsbkrcCy3L/9qNflpCd+/iNogYvKwcVNaxZRWH+n
I/Lvhc3WMpdhnel7qgVeEHHZu3+QKONb91GYy6VcDJoKsyO5aKrQATbEVD1VCBLSBhZqPRsdUm3T
yrsoQT72dGD8YDJJAqc4EgrcBx5ZpmdrQ57sDCnYagy4oYeVC4xRSYI+kDN/YJRjjte8XnTOROdV
ItN+IGrv666IKrPZudF+16xVMmphK3gm4zxJmfkppp2tHVXdUVQxIoaWGS6VuxhoPh124QEuosPv
oi5MjScsWXeTI42Gb+byZ8DF3ksjs5hv5SyErDalZNwHlaRMXKdXxsNxSBJC3m6QuyNhsvSmLjIV
Nb3yNetCgA4WV28USnHl/RM+BVkQ02epW9CGO3920TzBR7Rt0d7wNWcAJa3Z9G6ZJ8KHFLmLem10
sAoq90kliMSwaPttKmS8ZS6zbj4561ApCy2FyTMioG8NmPMqchVaLLyAWSCWXkOfK9JrE6QRflvx
fPnmpvrPws+firJ+gqioDRxI3SjAN15OmnWCM7Kz4fUPlmOYgTpyAJ8pD2iq/SWDVHtZ0obGJs7E
q7te9tS7Vxq//f/gd/R0+9OYKOJU9RE9G1lMV1/SzhLesDnHMFN0CrG1+Bfo/DKwtVkIiVLcfDvD
UL45getRJFieyTedIjT1OrvEs+Vd2dukKPEFOco4gNRBkwT2LwBKft5X8Vjqb6Ea5c94Gm79XZZo
+3Qg6V+XA/J8qD42fNuKRtXsVreAvQmWLJtjCsOOdldQpOb4AaEtBtY3a0os7UUa+usFQ2oUMmnw
GOamSScfo6k5ViqmCPRMPCXrASwmRP2dM22Bph2M49ut7dMmuJ/GLVotpyVVkBEase+iOYZx8i++
oX8PwVM2R4v76Pkd40vEczxdpowPwHb5Oxy2xXOnEYMgVw5Hh+VWrOhrlUmVATDgbj2fJf9GfErg
a8Ui+zsp3yI4L9op/5T9fdiqDLGr4dqoD/yxKIh13c7teBZUiTdkUUTNTmc/nbtmwa9LnmuaUZs+
E6ZZqw/dz7WwMUYBdLfth9oRFar0OJSuOi+dWO8KeVSakaa+n3QGlATLgMva5kyXW+B4em6Y2qtD
rShzlwkAxErKqRHPWGEnetts3X+nhbQoYQv4jR35KMkkhZjev3OtfncI3rjbYH7tWSd7kJweyFn/
IlznvdKl8cvOnpMHnzFqQQ+JPpHZsrzL/X8GiVABg0uEBJT3l3ltt7ifbcQHMDid48wQuLpgbgpn
Akoyye7OqqE+3XylBpc7xVNOntMSlMKk0pMMbPwHPJJt7Qn7NaZNMp5NAEWeY9LpuV/08l1GN+JS
Bl74qxjqbdW45LK7K97Xvfr/ubeEVvHTdW8RxH+jwx/j6twCKaGRBo7N4lHWEMeGT82AxtP46ga0
9g+E75o37wdmDM4vsrzmz/jzmPpiD3M5Mle8q6ZNpeMVB9/JPdfSAUc83+2UOApxKmJOdtThN4zI
PfOG+fAUOzLnYsGCWIFUxcK5BNsSCe6KTTwS3few6aBsut20T+igIyD48SO831u6IbNbKEGqhXGK
uQVv4aMozZvzOaQRnZlD71rDRnPeYAtlXICi66FZZfuwffCkz4HmKiN/TpiUhdkeNBYs6sqKG8sV
K1wgCyaDl71Nju5+BxTFy6KKq03jEAeNnYJuCLTwaiBhEcqgcWieZYanQloBtcZHU8e3xBeGTJM8
V1TfKCn2yGXFQojqhyfRwvGDAzR1Q76Cd2Z4WCb4eY33cTSWSjtSHPONoFWQOWWAt2GhZEyg1+cA
lHmpcmrmEukQ/7c3aiGjJNe5qDdwVdzfvQyJkAPifQM3K9PPbxZm2tjFFvh49fyAS/swvBOFZkVm
OtqqNXl8Rkzn7yfQGUXm2OApPonkfChzGanTFw5GNuoYmj0t6OgrmJhVtEsoQs4aQ2pNT46zHJF5
CUJzNTNustp4OShLSsxXmWSx/ctErxxLFbF6wvVOyQHrq3lsteq3xg/D2cAYaJDbQRWtyDqRo55u
OHVSOrUGMZRv563xLLyfLcDPZy4R1jwJp99avVCowVKwjd7BYRw3CBOtKjpbRQKAyrwp5BChT1Ys
xbm6Ga0De+LXUyKmAZklzRJT10x8CQHDSOys5SCzAWuqNkD9xnabJghg5EhjGCbXmT9ncendUbD0
TQlMkeFziNdtv3AXfw0JjqSmlnb8ro7kRlH93zfqLI0S6lWIT2amkaIu7iZYLenIJjhttO2TiloC
dABFG0WkBVL8NDCPcGmrb2sHLqE3FCkWm8tsD6XpSuaFjPyZZ+MXWaB4n0gn8R711e+7uBywFI7/
u/HVKlFH4eqLsRPm7/f5VQc4Y+te1+bPYgmTqgvGX+A1qV9ROS1vr0SbV18lxZp0JwfqR67U/S8i
raACWGo25gLKDi0eyRd7MimX5C5Cbtl1OMW9dksEaK+mquVMtHuLOhr74JPTqse3Q1CSA8I6T3pR
qP8Va7t9ywkxlU2YwiRoNYaiyQe0NAMH57OHJEfssL2iGxYXdsBmvfHr4qoNEnWEUQdkozOK0P4F
Mm7m2l2n1HV2B66c69TG9n9MTIGf2/u68lIZGIMj2rqGon7hmrjGHAbC+wqo5IEv12bbihyCHviY
37McMFi0opPZZXQtfSQXKRI1T/0ni4IiypwUYUCP7+4rsHWQVCrPzsoaW+cgRW9x5aGIxIsJjpS2
qrKMeSPacwh3IX4ESYfAcYocLrol2AG6vMnzyGwi8ysskGO26a6xRXb3Z8mdxpR5NxvFT3NGS1Xp
pn7/6JHGvUdfL+AFXG2Y0ZbnLKmL3mQkXPtLG8oCrKpXyXFMeoiDm0+qHa339moGn8osdAbzrRlY
H/SyUvey08HLeZnGpALj+HUoBAnMGpyaZBO2AxbHo/rtgc1YpDtK4mmMFo0DpTA7FNg2alBsYZzR
hyWjjpCyHMPUn8htIsXkLNFzE8POu264VuL6k0cV36ZaGtZcYk0UkYf/tTBm1nXcxrErXUu9XMBY
ryORy0ppOJv94ofXaixwsdoDUIVN2DgJ8fZntdLr+C4OnQ0K5xn/lgyyPFkuHout8OABotbmZRTS
fuir5Kj/ahFFPDmFezCFLAi0lE31K1V9TPXfymca/i6n6oizBh0to0idpNV8JzMeJodppQnv8I0D
giLaGzTnBcjvT+7Ten66KWoPs0r5uukgzeC6VFOdJTZuhiKzBhYdwvJqptShaS3Xjyw7NgbKz6jE
NT877m1o0ovNQu7OZZcyqrnHHhJDpfFjpgfs2nsCINQU4KRG2ZlqHY9QKDOBEky7ulTd2D3VRgpf
8cIqqoPdnEmyeTu7NBZ7C8wEbg+on84ANwT86iX9vZA+gYBBN2s76LDb7jahWd+ULTb+H5hSoIeZ
mMK4qktlR8J7ULIqNS7Hq0b/8yfTsfJHIIoNW+wC4eE5C+amUak3m5TJwYTOy9kh5TS7+Ba80Law
csKd14Pn4yQc/xAuX6Jxc6LVxpFZLh8dmg+XJgkOUlYyd7KOgNNdeXtW+uUQ2fWLrStc9+7gNWEJ
AjpZiNF1ReSO5v6mUaCcCnSwVjqwKuI3r0XDV///g5cO4vLsQ48AXxWHJAEajZo0d+IWfabRWEBm
l5LJc/bIyE72yBw43DtiDOY9JiIVo7chomN4MMWIViC9gMPEg/0oVP59YqSOru0MPbGglA53XR4R
m04o8tgKZGfsfayeF7GYUcTHIeNDtLYdAevVM9uFZePFzKsBEoMfggUWLiMSVQX643YHLCyFsgDR
VY2EfF4YT226IAKEaB7CjzsgcHc3CNWzs1qALvnphF2InlvaHdbBG34taVk7xdfHm+tUqZLoc3um
Av64p5IjjI4855QsH6m4su6mR9b/jE6+PWpTBt/wDe4zsm1V2DNZo+cC2ELX8oGgiYm3oSKpyZma
fgGDjRBEysc/ZX7ozyMq0AaWtKdmbY3B+jsHNrc9IZTLTx7FZujApe7VJAOiASKqy/1Fp/hvRmL6
94TIewJM2bapjg7USCRVx4f7v1LMEKeBCodhUvIjQh0YrvcokhRZf8wTZ9l5LLgYkYrlsWxAD93i
b5Xk6z8UoV4ErSzAW7xRPBGQrmKOdr4ILFEG1h6gjGeMVM5dfZI8h6//yrmQr2N3eI7QeqN5qGR5
4y0z9LrItR48SnRQ6kjlCgRv4tRLoqwIDKB9xEOxXZImJKksGYLle0OXC2+vYShfl21z/DSaPUH6
KGBz/cX9btr6Bn0piwgX9C0Y/VjB7VTDZrxIEtDiQ+c2vCi4sqEcPq3kBP4KjhyzIT530/5dYnvf
mu6j5m0xzKexC3wfDrXYU/6kez2DYaUP65LF2VroZzuWScp7PUxBmp2Avt0BHd75YjzIu16SuvRG
/Vt/aNLRL+wq5p1SUKoec+lCKlMFQ877e7ItCU4xzUJh8q/r8y5RwercboXyt45AKnH4HNbYtMps
udyStqTpGzpLr+w/JQK2yycBxCrujNXwmUbVSSb7M+PlynZXqsrz+AUjw0mrsVh53Ob1/mkfC8Ek
MRQhHHbaRL2rXQYL9UJMVVsuRljNCadqIVvU7IYz7LwtsTFAecR4/YVOjXhjgXN6I9hClluiKyXO
8eVfbpP34hkNkCKzRUn7xEnoKjWSl9Zsx1UJExjM6jp3GX8CywgE+EmP2Zy83M9utXJBwrYlKAk3
nJJJ0OyobdA5bKftGFxphxlQlgnI9/NYARMTuRG2/NUvsiGi5x/LiqBsJ+8TWoxbmHJS5XI1Bq/q
UQBEsEowhN/UlUjElQPaoONTamS8HcQWVRKRbw9W809r1XsYDteIwAcoVJOOBgmrsRkDEXHONzbv
eQzRta9DnpyT5YfcWoiY9NCapQO708SpJvTq/cz3GGK+zctmdGvLt7t9VcMFhyjoJoWX7q8hwf5d
h4cO3EWddcqqkhw+faLkDDKxVeCmlhCIwJ3r6GGj+Ntpvp06HXNXxvSbYCPmZMkwESJlHF6N8XRw
HTMjNuCfZ0tqJSwRyA9gpwJvYQUNZc/SbrDaQ3d5/0mblozxa7FUr/5BAs0f2/eh9+rcrT9rc2S0
oBWUs5eTiEgx8v1JIR/dgiiZK7SY2ZUYBq6ctJMjObyEgWme9P4mZzh8hXSJGoj8rIVC1QUQd7Hd
XRXpLe1Ddgu+8kZ48ykM1dL2qtn2xMICLnTvmTVNeVpJ0K5KQ9i/+kJdDGGoNRXJ5VwJqlHznyMd
dvlIW3EGVwDx1kKQM9AtNnEmEUBc/Oq4o6/CeyMLEK0rYmKxZpab2/LgO2B01XrlKeXFAJinkb90
RdELh8HV1fTFi2/0WIRO3UouWpLS7wftYv5OxvLEiwrIIF9UzKtI34uOxrmi98tNJzksmQLOQR/l
HNnK6TWNDlP2sZGKIuWC+HA6WLz5x5B3jJOq4rqit799aY7XCOLAQ1hMInMl1xptxzazfLystRyT
eq5rdnUggl1AvIUhCJBAMEcd3wrre1oSbdQQWe+danPrRBGWuxls44S8Ll0RlkIGARJItHEhnYHx
4PLqmtdfrTeLfV9+TQqdKSx3Yh0fJDN7CxB1D94DocqKtDlHHDsPxQ2rRk6R1wLLIDFD3rV0tMRU
kklwaCOQ96IQktPJgmg96Hs0ubDIhITJsKy+kjNAPPN1Uc8N9LLC+5HrzgBEuDIjCfzuYBDv9wCW
1Y9ZlCoik3ypAUzyBaSQa0h3sexUMTMyOTPN7XBXhf4nrH84ouYrB0gnjQj9AMXzly7/eAcO+NI4
P39FzKyqMXyE/vrfpMGZoBiIFuy6seCXxelYByO01OIbPhcl3354ZgeDonTZj5e2WlLcvSgN27uV
s2s93cF2ov+ekQJI82/WViR3i00jycwiqS3s2ayKGXYj8KZ+FsIfo/k/RWXYHtIAvK9UjPaJFwz2
T2aaMwydrrX33y0OJfmejL6RFIrMI0BBvHi9pAQfpVoWBBoyPVT7paZoKcICzTm170/AQWhcMAkB
EsBwXKqv+/pPm6KEEB+GizC0rp/kG8rVA7lhofdV9kOKwyuaC4RIFen/Tbcm1XKddJ0nJyB2pcUn
CJLhxbj7fdtcU2zj+E3bNcTDKwt4+M7h2E99in7OflHIG0uKayF85xmigdgIZ9Yv/SG1GRbBGpV0
meWUHbA1JxhYT3ENMXfJ4VfYfMrpOIXTuPg72RSzgTkXGA2S1MO36WzTaStoSp0Vn3XgFqWdyeBE
HCcEp+ux6QO+EsCYHX68/G6FL00nBWeFsLgBxZHjEEOixj3UWJWMF4Rk+W+IcOfcFUTewY9SNdA7
NCl4whFyp9WswEbm+j/4WDzfXf0p0SibX9kKRtVVctzOWpPSkTmMpyvl2AZSm4l83AXjpdmb6IYQ
KoCfmRXli6WWZaC4FYHgf/OVW1liaonckKURxfN1CleUBbL7/6OTDLlhxZJTGCazPBGQaX+YUDFM
fyrBgm4vFfvvgWMLjyiLY9XqO9dGem9CTCgZ4USID21O3SToC8FoEOR1Hw2gRKv52/+j0tlR4WFz
+ulQKaXRt6WZmbszy2LaJMZ8WM4fkdUbVTKZPEKzR+AvgOg5CynQfaYgdb9bkv1nhauxbl5n6R9R
p0dsRtN5z8pszlWDx1jkZOEyhFo2uvUgmvC28o0HOfwgFHlSNz4Feu4MwGryJ+OGZnJ9FH4Gqytz
BDpajh5uokGxcrxG23zQsSS+6DjjH7I8KLnivJr6VK80I0iyFigaIAXGnWwH5w4hoGzF+yLVT0Gn
qGcniEi0/lEsQ8BZ+yqD478WHCcgJ/7z8DLX0V6tVWiYMitHtvI6Yorg7d/ipSWL4w30pOlO6UjL
4+fcVvYE1mDoOi7nL8WkDXJBRMojpivotV5XUpgmKhSK61t5KQepycTWRicB1mccG8UfJNE+mk8t
Gn4pGj+limJ9FoacbJ0ePXDGSuZ2kOjXHZ0G2s4oWhhlBQW5STrgD0izEwQFZCxIWn1UKxWRhAZA
ksSpL2LG0r6uBydkLxtVNWIms9aDLQ6FnO5PKjOJSzTgGS7bHrju0NqH90YdKCngl8JoIFp96feo
AQMINj0wDkUVt3ixvu57739DHD5WtALDW2prLDDnzcsNhTyDjSKDC+Zl93YvyjTpG9xBvHR4Q0u9
2JYR6EZk+ISVwpL7nFCMsw/b087hH4KRQLfBnj4MBsRgEM/I+5S2LUV7ebtYkOpCELNJP3p5qUn6
FyFAfZJV+NKWaFDqskOEd0sNOubWdbPTVuV/KVZRK7z7HBEXmzOqKuRkQ1wE+1EEie2XoDRwu9Y1
gT/K4/zU/hMWPOIVDDVEnGDqhSsv1xv4yHyYNyLmitg4wmTd5ZAI45nPubsp4BNEiroORbZePVss
AdLNgrCLu3IlW/7jm0bOjo/5mY2cEfJv9NAFLOfz52mcudlGWZF5STd9t2w/CizXf7JF05zCuf2d
aQfBj/sG/V6I6Ff3Ws2W81ugqaU5YfhcbkRhw0hSUcCFnPhUgrpexrdVtBkoFQGxa3ZgJ4CDgxXV
l9h6Tn8epxslE96Oa4w3XENnEhgvUPYtEQ8cAGn/nIsVCHI2d4gVgTBDk+gCKlRnOIFY+rhwWLJ7
6spp9BxbZR692Vd8x8QDNhaSi90OB/lj1mycPg21dK1RUje+NyIahxZ4YHy0SDLCmbSV25/wbIY5
t27/1ojTJdFEVTHV9JgcaxO2PQNWSiaQS2K0hIl/yASun06k0jvQnKDxJnhxOM6ah6Y1OWOtZnfK
rQoS6qW9mt54dsXQCjhp6XVIYlrabd9A5RtI+Ln647xOspvVJgitO5IVEKuDqNbBFsyWonSmY6/K
O1C8bya17syNA8Lyb8OrkWEws3DflFlGyc6bW8UMwXYQfMM+CxTV5VmtWneW7XRgMEf6oGHJseoh
01UsbNDc//A6S2rULamxwNQqmDdiobfk/R2fBjamt6jFpUPkKhfjx6WK8QpE8gTluStXxUmoDSjW
SvLZElP7hq6BvVUPgBLuPWKRWCsXBtxLTdxbNd5FgvH9O7YC8VgVS5Y7/2r4i1pRuhEA/rlFtsWh
HB6WIHexx0I+mUEU85FRe7CUvc1TIBKsWoqWXFgF1AC8bIrL80jo+ueVQ4rHPcLty0+pyo7jqoHz
RLwwGEH+ClKW+nLaY3rG34tMhWbfq3t7KMzpLy+sNr4WJ6s8ZE4EBa/33iMaqSAQMO/HMpyL19Yt
wVWtk1Ha8lcXhNEa+Y9p6wC8NPQhBFBY+odIKdSWWfNf2XWhrHcVCu56Qvuuq6iMqfEqskxoLbfM
/MgqNJaWoTXCD1mhbGWRlmCitTHhILTxujfyoJV0DqP8IIQGsvW0VQojQM5dKpu1GI8Jj3LcP0s4
NTh4dGv+zntekcrTonHQRvEYfPdJ12AtCjtglilDkBxfHdFE3jEjIfP2nnlfNdxVWelnV5q2z8qq
hUP43VWC/xNk0xrzFW+9ywgqv1fwRTBduCE42tfnhng/Iu+3dj5AJU8M7LTMJVDHK5O9Gi0JtQfV
r8j3S1hNkvN8E5ono7h6FBV9xOj1bRG53vHEe5edq37/rKoGzkFwYudRBtsmh4kJra7hR9EQxx4j
37/GejflG6kDxY1f7xukK+uSeLfDiaAVSrPWvtOQkr3aLdKra4iO1XtSVlMocn2Ej9bsKHlMLJYh
PyW1f6ykET8n2+/s2/IhOm34xuOs+CWdKbCuGcOaSsD7jxQBCVVMfATZZweay3qjiMSjUbH9aJUp
IXabSuumd8YwdTYpU+71cvT4+KzufhjCfTlDXmDQEGskDlAr6Jtld/IiilkxK8uGBWaNSuWimHo4
oRkv97XJ1x8goFibUuxvV7jVErE8zkkMmRjV2+01X10+L3OEsfapVXchEpcnmgNiGo1eaeZzWHRP
0ruElNqqYCt8ISwupgYVFt/8WbtfR9Cv6OxGy2GGrEpzzj2STTLNcWb+LVF5/lHH2BIPAEtEP+eS
LHxEPLXymO23uJMpabGpO24W+bn8LtwgiAdnZJZcMM7ZMu5q3v9I+6B8Gnzjx8IdBnqkjAIrRDrB
BGA0nCvhc9EqsBwexICzWCQnr4HbT+zV3N/AFaLuM8/P0b84sTw3taCIJrqPvVbxIMBWueNFPlrG
FHwkp4lAdWT625545gxEaF2rIYipWbUhEI7rgIIZfrRQE2gBT4DO7EU3SSg4rdMndkBEBszTs/xx
LGMX8C+R6xd/t9mrpm5KerVEMTPA+0LomsTw8qlBw811AuGWjBEUZc4iaf5wBEQXH5MnR0JvSIjQ
7Bk+QWbksKGLnWX0dWZKRyZyq3drco1FeEovuHDsvA0SrYRiCfqC9om/5jxPZB5HILamQweCWWHa
xLJX02k0JfQGqr+LcaVmYmwRx1+oAjy/zBp8L2SHS3WaeyTUTg4Vy6FoElk5Mu+C/fahp50Bo10D
8hGN0OWztGzOB0xJplrowfgbd7z3JpEjYb2ApEmDQHcu+hBjbo7Di8TSgxLUBAkIfOyUcUD2uO/c
5QDgi8hqT1c/+cGv78aueJRjqtUrd2VmN0g7zjTcWWVScNL2PNfY9Z2oypEyaEaiVFJzxFNv8ZiS
wy7uLdz9G5K+lQ3Jyg5NUmsujYwEAURWRqAX3CVb+PMeAAd8MceQnghdb961JPIgWCL0BekZ421y
uJQUV1pkwxkA6mdKVzlrGQTmfXoThR++4hazKqA9Qv05DvP6WPk4zLgepDV8X475QOz/AOZDFdhx
ShUfPLfcZUBpVJD29e0Cht4eA3tnRFj2d/Y7+axXrCBgHHxFSLWDPkUv1BlI+yrRbd4OYsaGafgw
R+zOr845uOYJINQ72mBeQgnzW51i6KNa0U3yvMZdeAMUwO+lVOSXVXzMBEKV1JLLsrgD1+b5Snvu
NWas3MQzLju3ItSGWEwMyw5ojYVqCdK2bE68wYk8DDLFiyM8+5y+H/aWbD6xnJ4qUGBXvywoLNPa
ZCZ4qY8nFwNWTET3ge1yJbpd7jI/tFk0pJ6ckWZdhECr3Z7bZYvnGHRsInvyLVU4VCdeJh3pMMEw
gIrXhLQqOET0BdB6f3FEUlwQuaA6rx5AS0+mixlqwb2nKz7ndkyu1WvkbJWky2uzNR9m25clZR3E
2npEd7xhAyfiBXMMyKAllbno//TBH5vqhI8jJAEaYaD6AWPdRZgt6ZkqtRT0hL2r0nIJlXzyRTnM
PSEzTKKagKqui+R0oTw9WYd9n8SQLE9PyznfaHFOxdZOGMCNu3aM51XwhcNd1HfSbukGiEwBc/tl
otl1VAGMD8QtQni/lUd5lylwBXdtyFAQNCaGi07KBNcyiNFoMqy9+Y/xGmVH7CHOJ/xf5PqLVnTa
GiZv5mn98hc7xqUUZl441O8l9CHChjmFTyDvflieqxMoY3q+aeEXqmZOpEcaoa4xuXAD/wWpCRuU
1+5eFbBV3xDA4OHzSj9VHCStznX1HqBBdomq6gbI3kKFfLuJRwgF/aF/Ia5PY8EXNcqMZ0dj4+gu
uuRNIRUqOaDidvG9qPEBSub+Wg+HT3lMt5sqJZWhzMtFDqrxVZLVDTgFjaCCcwf8zsUVhTXzvX7b
6sT6wW+Ez95M75q8NlQS7F8bg8fLSUEHkqadmK83h4Am6eqUUhtJIISw+awXkkAjgR3xmwc8QSFo
oANb9YftYoSvf4vMDDnA8JorRaBeQuRe5PtLwhFKzEjDcjmg+g3sr0RUWUtxFBU0p5492GTieKT5
ftrnrtDOVqD/HZp8rts4/S4RSZ7cWzKPib9Ll8ffZh5wC11tyHkXEc36Exr6AiGKwOYethKEHip7
fUqeUku8c4vrKFpzNvCozEORTF0XJ5QKOU1M7/56ujBJXnnT/gN934NQSY/8lZSBsfcumYSklsuh
SSOSF5vS5B06SUi5ozAdInKmeN/pQadwOleNT5sWgIf3s6hinhcPVhgXKKlwhdrp36nXWZuwC6bg
+rJIt0Zo+4kDQL+chyEd8sqi6/OdnBTztOHQZWG73XbfOR4gOw20pbT43BEhF7h+T09kEj6ajC9j
2HSP3Et+0SjkPULiAXGkuMhNrnP0ddUuj2EjhYRqtyVRtvu0bsOlogXrFwoaRaOIGTbrPZMjNIGt
9kwza6fpfgN7aDwbfAAbjuNg2AWHagsRZtpnSDn/JP9O7cgE3/p6wiqhFJrNghExseiNZRfhlvjK
yZXv8/PYEeHT2ZHZA2/W2Fcr7U+pYnOyxDYJhZLXJQNaKPogg8mZkqCgX7f3ZGD+2bCQdp7/+/HM
X33e4q1GqjV2lasB6hvCBHA1NgS5Z12I2842aXTFQtYJoXK4As/PFjq0JxyGLX1hUTwhhZohlo1x
PMkRVZ1DjXB4iot00jaNFg20J5PVSJG2vShQlswfaay3royaejFKNTyTczo2Iu3fT9gowohW64QB
pccAroEBLp2+bl9XFobxhJcuq8qbmcI/6aOeJcTRYh+MOwjtNkfKq63TMUgssO+glFWopd/3f+Un
45JNjnNUbjgqlPzV4U8ARKO0r+OzmO3I5gNxBd50az1cTugSqEP+qAJpRYZLng/5nBxXkEtO0mth
dxGJrLkX2RxraT8rMErUb8qqaKhAXPdljG+msT/4r8PDl69IvJ+tFKai5kW1fr6ALcO7tUp0oe5R
XB8r78e9ghsaPRKgBCecdGPJpNOdHyhdLWAaaEa0PoGGxDw6ZXeQPD2F2VzKx6RCw/W8cX8UFOrn
1VX1zdIBrNDj1GHK8bQLy/uQ1ehS3pfhbfYyu5h6mrZcu8wQwhavxPDEGE50RBAABrVHieavOED+
busu7OF6fcgbxX9kFKVZo8MPSZs7T8ffc/X3uCZnFaXZyv4gg+HXB0zKRak4ICshC9WlZT2cQ4Lk
2pSbGedYCw8OPPKpDNZdSUYldnwD2iBwvf+btAGS10zPiLGyzGKbiVwvkh1fi4PlSiGY6eb9Q0MD
OWfo9TgSJEgrZxyCODfpswPsgRpGVq3utAA/5ICFmFfO/AlNc5eqqCVctDePFcoMHdetH5SQWFnn
0jdOumcM8ULTnCp6Wr1qZZwA9O1L37SAUZezNrpClUWmrNoVLfwz2Sup7nkAZA0AtefiIfyDwE6I
G4IuMPOb1m5jfqkZbE/TdkvcDpI5qcyiyvfewVytBxKoVBbnZkrnCA9PY4fB05EOm8saIDbT3opA
gVx9p/fExqGOVFABu4HE6e4cBXhyU1hdBniVP6yfjbzEKhHq4hT8AONGluquu5dXj38zGP2LK6Sm
Y2DrptERHbqyT6IT34S1KtEGu54YdeuiPHTm3ijBSQ12bMqUWFmenhY7FDGcPg7GGyDqdj9DBWXX
5RbW6QrkQqpEcE+gIotnviN4/uFdA14rsPqZN3yQtY+V/er3Q0mBUmDaM5mtCQqynAQJdcnBW82j
RWtg2GYo+FChqE0eS/0DFQJ+IG5mwgABwwn56ns5GBpPM6UQeapYgcSO+7M7fKmoqiVgR9zxnQp0
YNyBg2ysqk7CcmzyKklsbKvRBztjIrDSFwskBXD8h7hGcNjdSUdo/CDXMaRi/UJ3UosZ5SM00aIb
NHSHWjxtDy0M2DcvfuQtRUvFCamtbX8L+OhiWMIjC2xU6riZ7yBp/jAFMHzkO+orgx2a2TGZBeEz
zIyG5sh26aSCOE/h3fLRbdX4LnnGHtFWMgzawaL46mqzj5Itr28zKhnBtFjFbcmWwavk6Yeqyty9
5gXRRt3wVRSTwOkxTY4zXG8rtqy1TvfTx3fiVlwyzyh3xbdG33Ec2EGA6zFCocbURjNJ0SNA/+5l
9jZsmPtqZ6RnmRea300yZk5J+O/B9KpeDoApHAMKjhnqNDoeLfiAxYWTZ0J7UawFuDJXNAwVjorG
viP7KVQdCr8KgCIr8dgED/pLtut08U1FLrgs18fq3gZQAOfEQnIbrcBOIYx4BhlVbULDgzjCTbQi
o0zIzlcDqPzVL0+b4JDw9BF2pyUdi0KQ+BZfHj4Ei446auXVN6LXRYDIASgRw1fINnrFwGZ20nhI
Za6vqvcyNmhj9hwiOo6V3bMmBoF93eVEPWtEOmkicLkClzsPk6jXNYWc/FKboQ3Yr5OUBoNf+W+L
WFOu3oNC8R5aFSIHILnvcOWbfztmyb+sHMroYWjOAknhB6lWxZx6fCn5WKMPWplXmLqA1tX268jX
sFmN0d0Em6gtxLN/KHij80f15Yxf8ZU+GiWHZCYjHm7Hq+JZFKSfTldsJMnigoht8iJ7HnhFXvMO
LZ4kNOk3UeAvcDckJT6uMlUhzzQA4EwmxGD6EjSk/PiPSa7+4vzikIwX1eGoSMPtKtOzLRPcEuOT
QUz53nhaaTQlZCrMH/PkJtzqI3WSBcb7divxcQ4bLtQsIV/duUuaQtRhp/Gvrcyx1s1s9uwsWR0j
DgH9gFSXra5Y217AqoGz6uKiK1GdVhVX4T2XdxVUQwJb1mZC4YmKPYwjeLYUv+exWe+KcjGA0rQs
FsDgDEuLoIu495sKSh1qE7ztR7qqZnXTG4LlglszqWUFxLD++55k6OFoDvAymKr+9mIbA/1YbXMy
F/SsgiZSSVyTxU+Bqg3xW/1h/0y9Hllcyf7XHyfxEbHXOzdCGuu4azmMuffgXWvABsQrGnHKPG3f
GNdMmqieLUp2Hh2sZJ7QM9E4Oi6dfKNKOqlePbDTw643XKcIM+1vvWNMszjNeLQ4mVILDciWL0Sz
3eoN34eOW3UTAGdpi9zMz06X+LWpVPxai11qxf7i9+ONg7Q/LfGkQSMiAZ47ipY4+ylwt4Oh62oD
VRMk4jAfEiAX57UnKBUeutf3mjOkS2MpPnvWQSjUc7QToY7wa4cHUMe/j1xmrQX8xTzr2NfQTgZe
NM0zuXHOj47xSAlzcOBR0wXiMDIj8aGXZJGegWtcZKUzJnMpOIINGY7p2y7qWrdxzne2DU9Zl3VG
z+NLEHRj5zZHi4sBYjyU+ypwOO0fqjYkJ4Q3hX5zkz1azZ9Nkm7qN8bM9fHDQd8QsrIuebdcj9wL
n7oUSpo2Na9+L/3oJESi7JoyA+jyp1GlTSeNB4/ywP7H4t0AXgnQ3hG7HouglGqwToDwqn3gtQHn
m9pLjoe8ZEbhjZ8HPLPDXcefUNn+L61sjxgRFgn/VC/se//O7GmOh+5CUycHpnvJqMs8A/GrAtUn
ysHp19++1kRtPNCNnqjOlXRxld7Pdp3DhHYE1aladhk5aSdCtCTN9ykXF4dTHj6e9fN/Nz7SvVV+
+fbbWEQhH8Dlzl44b4YXQtRQ28fxDZTrHfVCeYX+8egPhbPQVTAt0mOe1c2u1Hv2Th1N1B4rmq8N
g5109YQIk8xE9Y/5zZJmr5HYevsTWQOUifRV6lLqu2BnhYUvZavGObfF/fvNU01S2ilxGVFn+PJA
04hOUqeF2zYRTLIio1rO1ahfztejtwj25ZP+QugoXUmK3mxNCvzz6hD6xI/ysAFFX1pPK75rpA4e
yftWZrcmvSDEPxdITD44SJGLNZr9t74ZX31lKyeCBz6KD0kXDHlSLiIPqh7seKjek3zBsAOXPSwW
NlVIY5KJt5RG/ky+pSTyC4Cbk5+g+09BSJcldB7Is22hRkOaKuAwmej5Fc4CIl6vvg1VN05T45Dq
8wUXYyxKw9Tv0SNNelyvY7BflYkb625S8Sk7+95pXfTB4IhilCNcnpEVNHcpULdqVwSeqy4CnEn9
K7fhG30M/ly/7NQMSHgEhp1QOWQWK6zMAmgeWubKUXWSM+4YLzEgsQoXoTt/0Mefa0DcOjmIg63D
ZRU8eCulXvCpJ4KPq20NmGGhoPjsDB+MfXAtjErNTOhDZJIg/B6L5AF/gbXTpBnP8xZltfvJXxKv
qpv+vdNU7BWjVXHdnw894AZf07RE7Fa51AQB6wFIYPNxMDBkBBIcmRVVPQlDE2gcpyyvLdW1PvRb
wsYRziFFAPwcTXjRrRqa8r+KIELFCa6jLeGTyVeYtgPuFX8CN1RHXxoB+RYDsgPwhoLo3EFY8qpQ
wFCSOFk4vit7dMdu+Pdt/2W2YYsXA/i86lDbB0ecZhEE7gR+Z/4t26NNvsDd8eOQTl0TSfzjZslE
yIsOLrzbVXXhv4Vcj9UdLKmvceeUPEQPz4JXIGG8QeNh8960gAXyNko2BGjNXjdg+kRZVJRGKJLY
oSov2LPXYeVnME+0FFDPAFTlZ9gRl+hGJ9mDiazUcMfpe5aZPcrD9+HQN855l5w4YinUqQvWqh5Z
J8ZXWIBihBc563aAOT+8eItcFnU81JrIwVM7YRLhMQCEo4F1FsueK1rv7pA0zg6OZrIW4gt+/KZ0
nUFuUBQBYi/+GSxJbZ0NNpnIto/TpwkCVMeFK4CO39El0wQC56yrp2unMdQ7H2L+zdXFMHL2vP6W
Jq1YHKbuy+ErgQC+dQqyHTwIBczbKEfJV1TSkbtX4lbR/bpP9wX1SNRQezXlh8tXMEU2tVos9Pc6
FqRXkiViQLmZAiQj74VcmBxy+6TIaHE8lpOKw6TlCKcKPt+UakDO2WX7bWxoKlM2H2iUHWu2Npyu
wcfQ2F+2oSROHRD0VuHYtNBweMNHizBE5TNhtSj+op96qczIUGxYteZ8ihpxb49BpyKhijL0p86z
tOwcwYD3jDX7anCZMe8KEJ4T6QjXHdR7WMq/LRmGCYcdf8jt6EjUbPzVD5wBApowlpy2wLwBgmfu
F92vrxj7WCt+PcOu/ZYzUL6Hmej2slPj6g0Wh20dZYxPlXfMJrwpEfpNU3iEo+65A2l/8OkThTy5
CY0/v0iV7BkEa4/UtNs8yTTnTTKvdU/VZc5TASubE9+UytlJDBXVNBYTk5oHZnocowC/8meM+HaD
vrWbXpTNnMHS1NJ35LW2mnHDTY2eU9+NMgAGyAVRCEXEeB6tvPXTi0WlSZcDg0WSuOrZth/+K7HV
Srqi571lEzk7awdDsdredgN2nwlS/pAL3+H1Vz23ylKOwswPmYyr7SF1jP5wzrsUNGwN6mPj7g+t
0QgXnJq5HCvnMUE5aRhwDrqNdwByqmH+KSB72JAcs+BhTx6nPCdSAW0fibrmw54IyE0Nt6oX2Jfw
50GUXYv2M304E2EbQa3/NzYnVkMkl6V+1wz15e/KOR8vHozXjn3zgdHVAlRTOkpu2ilMfYpGSbXD
VPQHt67Z5mCVbY2kZ1tImaH0UWH44AfANhtQ+hjtlxfy0+YWIepHck3RxZqR3vAdyyH4YuCky7SP
DzM6T8AXZrl8+eZ/Y6ccCmuREA1LuaOoZz4dWkmPcF0gKayFuxCg2mXkqYdjXajfSi4zi/VMd1Li
7y4LZnwsV4fbpf6bmvqXEE5QVYZfihAzNwpzr8dE7MUD1mSA/ByAK5d0im/8+GFLY7oVn/xYykcO
noviU8fJR+p5uKKG68GjbcavRcx4nRvlngy0cMh78SwPv66Qtm1zU4tfBu/caGNnrrybToG7tqoB
VkDsrnfjn5J6E/CC+lSxJ7pRUb+RcxASAMWOsen8vqOgYCi0aQ7R0iC2ti9VZMEfurva1PwH/yZr
WL3284iHabIyMpsOdW9F6hfX7RClA4CHXCE7tGsnuPgk9UHpZ73AxK0pjtlyhdxOyoqvBuiDtiVG
bjhszbWN2JgthibQ6SmCylkuU8rhjQcHGJZVFEeDrsWztQAvoiNHdYlTU1JiKau4cDA49Nl9LC/n
2/rapZgNQp8+KkrQccwj+bkDkfqVlc5s87DHIIpqsNQcDk5XlZzSp8bNO1EJM3mr9YSFDriJw5dQ
cxzn8m0FE0/+hQadfAlKnkMRHdOdCyuDoK6qJjfCt+qP1CmE1jDqAo8C/AhO/ejQTlRbl+3B1ewA
nC82uEZrriSGUuo/LDZi9DKtNwvT1/L4wEXXpP7JLQsacUlpubP1buupEGUqWK4PnjTwxLlE3/6A
gmitjFDjsh/ubnVGgAx4IAZ/G1MAL/6lK/nECupX0seEuZKys6LRHvtke+vKqUfo3BqfK5Pzhu/b
ehIuVbqNZFuU0cfyxETtBupOiUwhW4FHJ16r/N5G+HxgdCzfv8Q+gDS/rxT1/n0MxeK93Afdz8jy
UOhl3MJ9RB962GandLAKjR3ELb3pPPFhNNjc6AOYKo/ukIYL9fD0fQaXCinQmsSGXcdNkKo29h32
vupEx+ePGzzMvrWouOLQM7o0i2FsTlhF+FXB+cmHcvRbeOPPPmwcrAEujWd50Cr/5kAfgHRAGJwr
G4ZkPiajXwIfu9RloKJovjGB5zGHMD4A0AQzlo+osEtHvvaoHNMDuiP5UqvKpcPA+DRmb9wKX4U1
1KhM9owps9l5hm3kJFoEVrixEWbqaaaQ6cISKTF5MXlF5re2p0ymaVRij8KyNKGcPxNmn0VtQ2CT
X6jnETFqDGJUqNbZFD2qoFV1+d70HuM5vW8i75AUgOhH29ohBX0TxPmhHjQQLfgHIQN1IeVg3+Wb
eIgO2Hcs4Sx3tyY+QU8ox0f8SCGE04cltc2gIdj34IHrqAK/GZva5ljw7NklKl5wmnFa4FPWXQuD
usqgNr7bnTwG5HyMgiGoNGvk6UHbWM5g/JvWicHIP1GR4wwQQn7cuxg7xIBqCjjGmoR7JmFpaddX
jCvezvGcus8G56SsSlDyOh/Qcq1NuI9Jn4zZfPekab9KzIWi5+/YXd7m2CakouYQ2WzXPNpt+e/u
DGSzKIoup4D2Atl4kNvwc6QXZC46AOWV16HGkDWeCQc3Xl4rElwwbi6Zc/BB+j8EFrBUKj4S/SqR
hwfJEAcMLqQjQNKwyW+RbcHqC4yMvCQr26pB71gmTDrCKIWbapYweP680AIUPmURoQRSvJMsPdFO
fmWOHz4eGS229LZ9xB98I9KVLlUPCI2j2GAthTc2KFrtnQPQp9MxzN3SgWqzb9HUnFVjHjaPNhXM
ZK7piTPfZLyMY/FVKAlNBshgW3Lk3ssDCukAIq3G5f9X1aFRmtqykgu5hvRO7rq384kQiq0NpaiP
UUP44EhWeeWOdAxvp9u8XcXXFBKgeBfGK8pkFQ7HkDvspV0KgVtByhzpEEtNF2HjbLJ9rLVVb1+/
kH8B7FHLQl2f4v/6yDIa8P+WGxrBqXBmz57n0YodE5jG15ihvoxC5IFhN8+iaCAJhWXhvmWac/l0
VpZBlrhdCPRj2NNvpPmVbNckCQaITpe0i22b6b6paRjIW9T5drN9x18ZfCIkZwaWZPdMSJNq3e8T
9NFlh+yzQzlWEBYhjh9u+m0nAuw5qR9JgrChT3GcwfNg+hC1pJ+RhUneC4J49OQPJHv6yXFelTRc
Zrd9aSoTUMgBp6SYe5OCVK4FIlH3Vsjb2fRQACkD5YYPtcW+apPs/PlN3y/WJcXPxu2aN3o17Snc
FXNPDHhzrwpAPfR2wmhUN2MVFO/M5OIQH1fkoqocAMIytFRN4wDWO8gU6MVLWB1og+vKT1GhgltG
/g8ljtW+adQR9XIayqu6AGQF/zAIqKdcBVydJObpBEpUqtnoE9HfsfddmvGmEqzE1J5E8u6vgGYo
/BfbDJajz8RD4/5BJti8jhboQDnWSJp+7Xgr2bjA1P3Zlb8HdvR4W/ool0/BA6CR0uRGYC4ahZXB
45fyJo5z0o9CoTxiXYWv9lPxF8aQ+EYFFAHMquSEY2CirbXRqn3QJiH8VqtfxItNA8eCC9m9DUDP
yR/6m9WDBK24xAnQfRIFyZHGdWyenKILrkY5Ulv2vqIgyto96rYWUBVirWp8MWQsSYkVeKBTmrjp
eAXKBTmhaOeKe82MSE/QSJ2RQIKnqob1crEmUFD5oVriFTDCQudrnNkywrUxdLwK31muO8VAuLka
jFeaFxcrSto4wDrlci0coRKcs+xE2erLxCFSxTT9fbYDl9zt1cH9LqTijoSdUVhBpLJTr7fOsD9A
jEGlLl7PX1WJAJlh7g+tE+NqQadIbOPl+skFghL5UuTIYVVXb42i4+HDDhS8AqWnArc0uz7OYyHQ
A+V0UOyL4ZfDlkT58PMeNiGFhmoE5jCq5gXNsJp5iVYfJBQ3dyLufpMef97Ik3BBFicwqop6GfQm
m8aVZ0PvkiAJFB7JFI0NPbN8v6goi0QpKkOD3I880IMSyboo83cPhcjYSJXhiA00s2mqrvOA4HuM
zerOgtZ+W1LTj0RfFulKhhfoX+szb6Y8MGzl60P+cK+EcERRQg7qvHod/Dlrb4EMK59qtwHQjymJ
IKf6AnxbRbmz4WFi7HHd63kVmYBdQdQ6XqnZbQs4HpMmG/vfmEvK1w6405ZrErzvANZouKa4u0K/
X0pFM8jNtO6ffRW6pGka/umB54f3WCmD4h/YtIQvPgtMtx2XvSUFhTCsTWERq1MkxgbV/DXd5sAI
mTBEihb0QiBSbBd+OLomyRUX2fnCPkxPsNBn28ndVDtWth8PlmICLaEpLmF8cIRqW1231bGmoFN2
RRpJ6q6s1scxf5C1UZtJ1VmLOyY6tcdRr0cUsPSTdfIVK3rhH9S4jWlQKGZpzi+BF7wK/1u8egzu
DQ9aFiEPFy09EqMwe+GUflPLwI78DHuo+pPty3q/s1h7noHdYsmahwrisHQfe2jFIF1Nif3JmRB/
QYIhS1kjhnFsHu20Xz7rztO8gkjbABpeaNIAHlRbnXUdIFZwVjTfiedRfYb6t5A64TxxDTXispgo
FaKNKaaBBemgkW3QF3uBBKQLf+s34ZHwnXJpC4uLtVHhmfsWT8P2UKbA29sEnmvQSM4NzwdgZa15
y7I6H4HKEwMY1NVTeU+y+skSb2oWlwQnA4AU9jKgjT8cqOO+yjsVAZ4A5dg/YXzba27+b9kr9sO4
S2v/RM8+ebrLPw+5yOJXE5vBgX/okJsqyEWBWOeycgL/uUPp2pfASgWgtctSPxsi+cUldJs1nt3Y
W6pAliUueFExyHD1MwRkpogwpGt4rlxGkZD5MN8gsKjYVEakkNNkRDZ2dk3+guCnl7ikCoTS7oLF
z1Qux28fk66RYMm7eZFxoGjM/nfpqP02AqnlacTXhHpCP1wZxXkNXTlY+uUpmJdHDZJL601wdivy
F6W0oNCv2AzuguUvCawEBiacK5tbL/MKqNfEMpSnxnG3x9RgT29/E/4nXiYqOP3AD27EXR60rtzk
9e0wIovtuS3lhUMYRoNxxjVymjO13V0o7UNhmWBIlERAaxprR+8hRI2koy7EzLPPaWtEBglO3wPR
6ijN4mk9gKkWLb8oJ4cn3mk7F54Q2mimOteC9xbPKIfwlT5cuMTcCBD/fo26PmsLcsmVIuDdhD/T
WF32sWQFfWQg1i6Y07LVhrWI32QmDesf5EU5KiK6uBPkyVmX55ZztpeP41nbxMfBtd++B9LaaSHy
KPJoZaNE0+MS97R+woJtmfYK1EYC8H1J2HXSGdRctuYrsotz63nkMBd/e15XQq+UeveSemg+04C/
CJPKku4ftXMUBvIN2Ed3fRXvPOuXsNK4KHvI4iekE/G2tNay9P2cVTdeOKuK3Xm+vh2AVq7UQOHX
Xdlhgm6XxPTEbPVGTtAVp+TXiBGKVRNa2zOSyLcE5pSuMSXinng8/ixhDGTbfmxPARE6vmMeY/QZ
K7aNlH8KsFRl2NIEscny+b7y95BupHxTmCACed4J1HCv57Dz/JsPIG1peNfvYeOzOn359VncytfF
6rZGKb7DQD87hC7Ln+CK2RyzURKpzdpLPeuqq4gNal3/BQ++PcROmyeTFl5Br7rv43R5ebA+RR/E
eRMbfMhrOVewhBe4nwANolhoCaUi7OS0CJVpjiTRQtWJVEFY4gAHEcO4+w3P0TXF7Q2LT93aIDlc
1tyftXLopPO/nJWDjRge3IilZQseRBDChUsiOEXWHL419SGC+f4KheVhgLlGy7RLTTsZiJxHiQoT
UJmpqhg7Jmq++avqJuA/WeG5r2/ozK/IKNiPr6RyyFR8uRGXFAAhXRuNeg342tNerK3CrZCCZgPL
M70Z2SWzngTyj+/F+gq8aefOsj9LyST1VU8C1/Fg7NDQTS1cQ+o4RniQtnhbC3nR/5+Jt/3TXuS6
SOgFLv4CMDdrFKla5lhyJd6jTLb4kVKAyzcD6mxEIT+nh4WefuHOqEyKBDeg+S6qD5YIvQvM3ixB
N2JjhpDQY2UheGPauVDajH+Ve0JppZ4EymcrTBUEilOUxeTNv7papHuMuK94wUxfsCNnvndMNWzG
pHpTSP5CKdtAAFmNqAP2668jpC83uR7ySD4OJAaK0pLX22xxr1lBGpYqFkEPxK4+VitHI/p00AZY
eXZxG1qbSgqQQ0wixe2HS4Sli+sXW78zofsSSyRkiP4P4WviRN+EKhLWjWaJC5zbbNinkuvDsfy4
c/4juJUIJQ4VnVci0OLZA1lgM+EKH8OMQ95hAGnVy7W3qlhWI1vfs1O7bc4GlEAejxw5H0LzPr1m
a8j2cCCDXlYrD5P4sFLVA/QjkVfPcqgZNtUk5Tp+aFz6lywFGBVfS1vu0EVQ/vQeCfPbs4Zzkdql
yu/psTaKSb+QMokldf8No8CO4s8sIysPcf7bjNxYaw42QfqS08TvsE3VpvdH8ydLA/m+Ya1qf1Rg
woJ7BFAclGYvsWTBzMQNRXM2oD7a0cgpP8Hi+mafGB7RVdWSHV/N6Gr6p+/qYPLtVS7faOIvWPNu
zY4nrea0N9LEgbIvsc76cVbEPrvbMfaptskx6qSvGj1o/w0cK2rKWIxLF3IZTEqsfY09JV/Ilp2q
UHA8tycJBwlknhzCyHbnDj1xWd3Cn0iAjeZSHDj4Ot5vSMz9k3YN1gY3p8B4ucExZGtoSSkUmmnV
LfwLVIBCOtDkzo/GRqn2Ojt+MTRiqv2ECcJl1sfGBgzp15vtPBKJzjHCancjVRaLTl8KDdRCOUwN
bUWnB+wC2aEQvdbDHzWsPPtjMJjPWBSEOGGOvcjb7V2bOAb05yRPZf6kzBWAY3utpQb5BrCzeAPc
uLho8DDPNiXpyBO6CjcVhafORQYs4buKoKkANi2fcvse2JmuSRhBZugEHC+pIJ/xQKR6QWKD9z+I
3LDTWwF28A5PtqiOIxJDQBfxDUKWYNH4HLG8jzU5LX/rBgefZ3awxFm7OflZqCVkfD039PTNMgsk
DVmYun8pN+whc5wW1HDlCO3QNLG87e/PrJlCInvwnUgXGHGyjskoFBv9tSSqJz0VgHRIlNyFPQt5
7njx2of5YSB/72s0dkCztsQ614LYGhrLIL/cEgEzpltsXbaYbJ4GaIP7Z96do/EBWTPq+ms7/p+x
caPY9updMtP0JhO2ZDr62wBftMKqZ+d5tojILQgoCBYG3rc0bCXvCj8atg7To7RvRmNKWxQq9Sme
SAYWq3yAtjY0QV0sqwo84ORTAludKvMbBHM+4Uqb4Bh2AZiunB3U/2e6hoH4BrZZwg7KdxPQ4qne
4kZPdkDbsEecAhgNzqLd+xiIlgrI8Ad828MD9MtDjRnzANU8ydKVIF44n8NP6Gba4JY+G1MGz2MU
RMh4FkSse/tw5A+qTWs3grBBsUIFhInj1sGo8nsCupENurtbEIuNfjJ/wB2OxIQMk69g1iC5hvip
sFTkt6XRfDIO93rzxAhOv7p3LWTGtunw6Hqk/nNtUzrXIKfmdYghDjSzhfGlWrM/S19NZkgnAG5A
OIsD0bme8kbD7WMMfD+AxfxRjUsqfNjTggCu0HuNMRWY7suzKUkpNQEpdDGqJdek8JX0yY1LDaND
XfqT8x8pbmhuXlHWG0SZIs8eHwk3VMfpSSP+AaH3eS2WuhhzZhUWUd8KsnhBtpgMJ/LPOvOjD5MO
zhIgC7vcwExwk6j/RCitzsgNK8XICOOToY7P4s1aAw7Wyesw9cwLAHC3qB/DRCLfi8Yc8FQhGjIZ
qBF70yyLsG/ucKsFcc1MGkAVzWGsjGMVvH3fOnm3OiCMoJ3Rn9wZ9uL2DDsnzPZlJWBmxSFawDWA
BPH+Kd+zKm8FemsJlNz4GV24/SlKRHNgwHSOnzKtGu38Jr3aBs7po7TpV3e9geKq9WmR9F7NGhkw
f/ga/Sqn4Y6kS7cxP5sPT122zCN7DdKTk3kIQB9cCFTTAjE9VARGM3Hgg3xmKVqJdGQVF0j6L1N9
L9b6xDbo1cZLhmE3VA1SM+CTEPPNu1mcCJ5hGg/s0+dwEM8Y11c2aZReLWzDfgI92IqQcKUC/DFL
/a//nqesaV/pTbkaBW+ktUxdAgjAPMFfP70X92wMVOTf+UxlNn6H9wBqsG/BMMIyzeAP5PtfBc4t
WeUDcUbBLgugp2EKqIsaGjv6Kc+kW/An/6Pkdq2Ssm+CaZJNFtVHHv7gt+sC8BfrN2q5Jf8sBBcB
+WptcikqYurDtev2DPyMDZxVcpnHBfLsT4mvE3C8/mHJTp2yiMXqHX2S72KInKqDXL6TR4vU0958
rc4hwDtBhKSnGIY/ENUos6uz+xAbGyhdLItmiYnGfgLAzOYxrdJL6NrZcRWFJeBLiFyAz0So4a2G
P8JOBOVJVuYTPLefA7qmsAGJqYWoujQWXuBCZjjp+YfVJZNDoWITCOiAYlap9KPA20LwacUXuL5J
borOxALxE63wwgPeGvHe4CPOWY3x/DF63fGKcGVk8o4HQGZGKK8ET1pfQ5lH59ZNVUTvn8tigmce
6RnDj9YpPRWsvy9Fe9FWwtl6tbxDomEyBhW9ZUh2YlSMjmKs1TWKQk6SuMvx8EH4Faqj24togdBc
Dpy9ibo5DuCMb4/b/qhUszR7Ek3c0ZpboWHMgLUQMkAU0SXrZhTJwtN7ZkLubkw45IX6zc2/DzCU
88g0Zl8q4/qvtayfpvVxeyX4oExB2kHbSL39V7E8R9qyYsR4+La+AjtYSxAZSh2AuOzmscHJa6Ij
6rd5a4aw5l0Ee3ZMi3o4gj3pA0BHyeTLE4Dlu1kQs/jjI5hvLOwNiVpFaNHsCL+SaSfB9EwnEbWM
P2eBZmh3cSzaU2XaicXfkTt8vhhH4ZW39TyDsJGxzwXuPM9uzVFXhHh2aiwjvyX5fC2x0dmwTPyR
whOJLYrEiOwJnJej1IOWNICRzYKfTEVMUSzCJ5jTw8EV55+OIZJP5yjyfajASlj+7sbI/YCynmSX
LwEpuOCuYl3YERRd15s6Oa9E63czWEeAIV0LRzVfS+caVf4kTYOndyQsmQB2zUdlq1fre1kRr7AA
0p7qlkoyo1IEl+JAaEF0aEDhsLSnzNTZTQ39+fJk07z5SqmVxB02zY73RA/VEvq5+yNgq6DaFQBc
Vlye2tYWUyRdkYUGLKrL4k6yvDCa21B64tjEY1k2Iw13JwNkxG1rqK7rrozbChwnU189silmy/Ao
4A0T+ZSo3W0Ecq1SrzxfvCiCQ3vcv6jxsQTRDPF653HLojR2GpTaHqHTPbb3S18YfFtJtwIvBHJm
QxERjgS0qM0sBJcuvwtLWLX3t6uEH+FJzyguS6e1AH4jw1kf2BXGCDdhlHHXuFGHeGkVy3yZkDYZ
XU/ZVu+bUpvTBx447oA9IaK0Cya7Cn6kMN7kBzekQ9OuYqj39SpXX7Q+ZfFxHAWUXBgRMPzKHYFw
0+ILK3qo05fD7L5yMMQg49BsmvODL2anK6w/EcG1UnlVHQeqtG3MmdxvHeAlhTpWXmejSQ2aN7Dw
vZTh1Hx3mR44CqJ4vopomTdsboDxtfF2/Yh2Dj0nAjuqBpQzXGxXtDGbYrSnNDmIl8Z85Yqi63wl
okaiFfTFaLRURkI0rNKVuPgtbpHYRqVJ8H2T4tbFswgSTFvrntURp/IOUWNfpcOM2IOGLqSYn87Z
dc6DKBfFxr1PlcgO7bMziWH7IgKhDI2bd03NrKQhF60aJC3tqWBzPf+k28cq5aXnAXQQTX/dwDJr
8p9dDSTpImmj04UmaMZ5l0WZPZCSHza0+5g0gNr4wEXCKBLdGSM4q+3ML3K3F6OPQ+nPsGPaGn/6
BpEeA3NuM2pqjPsx5FP9XaBm5Q09a4VUk7BkgAA2DXk2uBQ89ML0/qf1ywnnzTvo1ICXNBDDJbmB
Xk+yxZ9Cb85xCsSCQrzyaEgyyOYpffO6GHpBgmdRhS7tUspCUIcsILo4ip+z4+PBZO3ZO3HWCOjn
ty6TXYP/jmcHQkRuTfnCJfmqHcyg7UHWI34RiyEK1U0+EOZovDHYt4HJ/Ck8BNbsiCYbbnwKIlMY
jsuL0AfrdenpNhrYEIjm5EbNnW8uXpZkdGOOzQfwWIVOBMUfmQ5K80VKRT6kcFAyBNh40OTCEZ+x
YO6OsmClYEga4WslizxmxN2ywEPvRE+sqmshOcF+UxCgxp/ejxLGqgi5+fuMrqN+eGgOjWpNwpXL
6uP43ZaaGhyrAR/I56GLAMvZWtEabRsovAon93N05jEZyAgUv3F8vTw6iweQCqJgGQuRMHOnGQ7+
9x3q68nDfAF4f84gO3efKPa+VAzK9HSvph6Y67cRJ3AKVZF5sTyC32906oYjDEy8YNSYvP5Zl0um
l/0PI+xViYv4vD3VXpfoKTEtPxbfSIne6ihX6jAvH8Uk577jhdIWobvaO+v5o2zOHhEXId2SRRib
4evdzSKK1d4Baq8vg6VjWgdzxTIcbKBEkp1muO4fhY1z0zN/zPc6KxgVwXbc74bYl6gHpxkvtv73
yuatLmtSEzhckQLNqnVrkeeRrWoQdudTvF3j2Y1iV7jj68wR9FD7MHN2bOsyjsHGXAZO0STKtFbV
LqBCExeZDuqwn7CQ+TXKGUwk0/+oD6O0mLVgieT6r6eubyiWW2ntGoS0sVI9WN+4uBoGwuKwyRA/
dk6HVdREG/BawmBtD8egveg5hOIK56Yr8WZrca8wEwERQ/gCr4HnFZK+dVYsZXpnBnIm0D7HAefG
EE2hRXVP61SzruT+2pYjOJufbk7v4Vwqphf1pq1slJR/6XGTpjjDKjtzeUwlTVz4xC3kT19Eamce
nLAbBRXnywFTK0smBHMZiBXobreixZA2vx7/p7DSvIWzvwBiffJrFVvCQ4aLsi0OuQZtq5wS3uzt
oeF0bVe10OUqaO5Y6F51b9zd40DnKAvOfKx+y7kXXY/ZViL2fdXWU8tgyaswQXvkrlGQX15gMKOu
4atXvfWUaShgs29FrNc0zwcGOHxUar6Oqj8W6CLcxg4UwY8Qi4hVCm9cDRoFzyWhf2XiSoXXWGJ2
miLC+fY7G5SwVhdTvdE7mgedKePqWkPD63jwxPKJtVct/tiITn5GWBsmp/7xLBIPWK18qnxW0rqw
NjY1jMkUPfSZQoa3mTDFaeRZteJJkcX6qEXUA9yORbmgG3OAn9D6N1lOWS0FiNOHFKYEwdOOiEQw
AC0kmyFG3pPP4LmNmF+dVUkiTJ0FjJgECZB5BjnTpybcAUsJ18Z8Kskn1FoH+ESLSaF1z04+jC4u
pfzV6pz3Y3QQ9EWP4+gAHrereK7/dqyQdZWllklHW8vAMGBG47yAo8BVDIm0Rx9kNhMOt+RSe9jU
q/Tni/PfYqKTsn9bi3yTAXYQ4K6fRBI+ayD3FLVJn8D4M79x5Rp936zi4C5SDOU6lhvQrXs71kHp
yaECmI8alRW1pC86EaJeSmQiAFwdvW7zhT5JHRYbg7OnztoRiS9TVLosRuvTLe+4PhLhQHhktOTY
j4kkIwWQsDWWBTcfJkdnf/9Z8a1YZJ0e+Jle6DHx5JnsnrGYff794C1rnJQf1ut3xsRLJGSgevkp
GKXpB38aZ1maedNyYNJ3ruC0wxh+ADpDBWkrWQ85YMl1SxOK7MkB8TpHLifKHJGU7IkTIorAsGc7
vXmJYVTP7JQZbCfwDoFNNS2k73TfEkPrgHjsL+mZOb9948BeA3gAGPeoOZHEYlXkAQbejiHIRqLc
rTxYCgcnKh3g0JhYIwrbcCbZccUsulJsZDJnA68n69Pexr4403cFtReqyYxJjC0mmA2nDQczA9Wm
3rkjPPAwEFKXgX3thYO688aJAiKpxg6kL7Yzs2HkoWjjnglVdUn3on7ZMo78HkQpLDYCbq7V1bF2
tzVwRzkLWGUSVuudbXFx/wwqfD2f2wHoWFeneDfWYVlv5YM/DYfIVsM5Pl4/FccedTx62NxX7Fvi
xw+Q2MKglUTRwHx/YLD8cNiYhJqvWA48qSxyQMtlIbHb/eOq65SMNlEseqcPw05c68I4wlH1AYfT
+2XXbGprVeaa5XGKcA0tg06ycbm4qCaoREQblReCSdYJb+VOCOK549hEzqn9kqrqSuhsPoiHYjk4
bJ1okToOZOKZdsVnX06GYjYI1hbfqdga/S1BRyig1mELzBwHCJmGOSGYBSyd7Qyxy8F8KlDQwkV1
lsMi4Y5KUjUy2CqA4KTkwQ1yjXkJkhtjZkVLDZ3xcUc4puik3rewxnKVGO7kuWjkKu6rsQlENO7M
xl3SIFJsS5ooLkFfN5avNFP3PcDadR4IyMTAMtVv2ojoEMhSrzgkxgboNhSy01XwQjGoMwEtJJLy
w61PdcJOvpNK+3/qfc80ji4PGv9xvARuXJhzNsUpEPqW42RMYcrGhmzJnP3rSmOMMUiqEiMtRWh4
A12vIFWxIGGHviSfL5t82T+XDFkAXYrPiBFjOyJ318ydDRT2CDs+ybcdk8bEnCMCQA7/apEwSf4V
flNEga6CUJyuFLFH9c9jVBEQxO5NiuK2yicK1qnfVmzhX9NNFPZnklH5vT1znAHjdMlY4yzhoiA6
JFoPih/mju18dgt9Fb68Izj6zJnuInScHKC4zO2sb/ECuDI8SWMiROAhiNMwZT8Ogtd0saXRZtHm
Ua8Q/eYloa7GYhnLWfL9XLl0xRNJeMbcA7MiAfz1cu2jwQtrB6d8ys49Bqep7gRmd6x1dvGIzb1v
tkd7TVTh4pxrdqC2YMrCZZYRMigLEbgaALXkSao/uFqTl9SmAUOTMb1zpFJ3ciIZ93PcemZUvOjX
ndLKs45dGpQ9MUAspP2QCxpr6wXUr6MQApsOhdI2QdPdLhFRcyVJKzHwlweVZOlJayUnfj5DoQRT
qqbWuS6FbP3sJkcVGwzYVpNkFIdHp+yx1nC3898A3gyEMpeiz1rnxEKA9IdFigX7puObrxKIohOC
KiQ1vmyIL/tvuXraAojhIXwrhvH2N3oI8BOnq0OLiBtBoRiv/yu9BSvZuQjipy3/zPU1Jdb2WxnL
pTtpV2GOoIwHeFpa9RAx6s2uz4Si7aNeQP3FgdgVEowYef6qVQllTIeZ1ip7U7W0AYeGFocNlvU0
/PRJPuVQA5F7VF9XDXAzZOktB1ZXSRF6ItwD5ckOCixYSmFTc3tYg/KiYZ7RGNfrpQhgHGq9IY/w
O6wsm7FNKwQL6o2tv73Mmf9JJ/RCe5cT3xegW+nbpdrxx/nQ0rlYoqvSmpQpPSX1vuiJFRd/pB/s
wHQGPkspqdDkLZmTtcQ9PDBfUQhKGNs/ZYxzAh4FMYRRD5h0auMloL+aAy2O2eIGLYeMv87T6w+h
M8AASpbZaVQtgFh80weK+YaOnt+/5h7vZjHZdGmpG4pEwPgdot4ZhZtafMdFlO2ph2R2TgwR7FfQ
1YgmgFK1f0pomGvqHfFbpUIqPRTckkM9mdlVzBje7KDQxSYuIcbj7FDINOjA9ZWLRsRcmGOAUuyx
edB9ph3EOJ/JiKe2YXaYnHfahj3UgqwNVMcCGFQOVNnRVGCXT/WM3QgRE8R31QsAGOEsFdO3zJ/0
pvNuoK/nzGvygx82G3oSuIug+afCpC6ZsjL4rzOAnn1NuIC9G+yN2bNHy2Gk/V/9ZiGC/ZhF8BHg
369GhRZCtGUjt2xQ7xwnKOpoowv9ZypIJ89SV4IYvMbHG0LydXpYiWo9oIAvE4P+Wao++a+CUVu5
ZsGpl5QASBvPZRVzEZETmz8mXZlUhvef2NL8U5OMe4NxmLPv/Ea2QMFab6QnGD7IKWaJmTl4gVtP
Z33nn04tP7XLIFVLCeTNrCgxzBuxUDeYW3gwqHQkKnXfmDLNLmQRqnohbtUs2zkdpiBJzgLsNRjv
C/5gtHhxWgSrhrhdKD0SrVbKWaCn1hfWAtgP06oVelLLHp2SMqBKpFxmNqgjG+WX18h1HRxiFgyV
8KZunOsf7T3uVL5wlw3T7zo2J3iseW3+MU1rCwW5tlQMAHCWimkK3mdsXWnlkAfk8wq2hLfKuQyL
U+DSZS66StTfi2h9YsoKd4KE8pSDSb9nAwfpgduihiWmd+HqmqvyFa/OuYRa3OEEIF72NAXZI9mn
mRqxU/BYPAzFWFOoqEHcbYoMltvWG6CJAUmTHMp/gbPszvPCx62kkfOP7BdYRJX3qbgeMHkVKqbs
NIaYU5i1Pn3a27sXFLBH9In+X7x5GPb9WRkIRi45F9iqvk8RUcvm0oUX65i2cWbYsogmn5bhEmKA
9b2ZWb21HJVktb0TYv5H4EgqF2+7qKplMxlRmZl8iaQQPSyiMe3Dumk6kBYCh3jagXngEnnqdW5U
jjD01FJ9vuOyoi2PROx532+vxurPRgUXXb8MGnz1dNWXSQBirNSBgdKilz6fd/TTNFbr2mUJX78Z
9jVrtnmjLl993G6rB5aGDlsBbf2V+gFCD5F2XVFFE6pvNtKh4WpdjfU8WDKiYCMUX3bAizQboyAS
Cdz/XJJVfg4cqXOVdjG40009xM3KEkq/8WsVs543xHkxAP+/GQ112TTjeE5Vhf7QkHba5TFX2yoJ
Ep4u9ZINyQ2uUkU9ioHH+x/ORzbf/iR7HATdEVmP4ZAasvwYid0l2x9OjJXOjcA7TSundOJrxFj4
qRn9eCKMtpk0WGhztdRdXeqY89XEiwJZ3DS7YkQ3Krvimy6nloMVNSb44uriO2a/mvWB6wcZW6BR
2aqWYdwe+yoxBYrugRnjKYCAEaujNjZfXIVAZK5euIAXTg78mcFsP+MkmXe5xXfABxf7zuUvLuG0
ULfGovrfA0iKPsa5pJAW71N9FtI76HDPbDY9sW3NQYvhPnR76eY5Jk+QQ2hltHlcEOeJWnFeWtcs
0ZBTlYgDUY9WEmMA/svtBDBoCQgF5XJ4c5Q8mCNh36msSFhtnaWymZAoeU+eI3DWz9YHAQA0D10d
MxQSAWIESlq9+L3HbdInQ0pmY+PNOWYNXC92EZTITSeit/xblnc/Q584NjBcJV6ACPElvIXKpikQ
3zGPRHbfxgggHKmUMorwHXA0ObtiTil78qw39t6FTEbaJi2dVS00pSlZUs3qHb2PEJhTRvuHQ2jo
XuQgxZjMN2/NKC0JO9sbMoZa0tCpFquAPD8waLYM3E2FZ+SdahKV3HTfVDtwKudhFgu0ulU6vbjz
2zt/uAx2L1v2kKIroQ2SP/dVdxJu/1VvTl+I/nDjPN5NGI9BaFXqE1jNtMvtSlzw73n0DowiO9Mp
3SGVZXs/d9ec2oqFwHFXFzCslujhWcM16AlIrZ5bGxOO+K8kARjzu4H5L3+k6rOXPIrxfxZzCrnq
0at99R9l9zg5eqbf9+kDShlX8CjmjoN28NGAOootT7A2bZ//QPFM754oV7ktmH1812DKzTvPlijN
tLM3evJ6f3y7sZ/InvfAmgKRTrX9MG0gthoz0OsLWr3hz8DVEZSu1MbdCuuINKgqeqfKJSvi94a2
daEk0TBcCAKqf+wqWuuuQreDdI+1X5R7XdXFJ1i0HlNP/iajN9yNreAlYyY0zyInKW13Dn/FKGby
wbUdDXv+5V8RBkh4rZrMvxpLKSiEUdovQQkg5j24pAAQvmDbzmUFcleQZwEnTs1+mJnZdNVWUool
qQ7xes/h1TKyya3jhSSDS0/DjZH7xSPoEDcyopovZrIvaARcj9f2JTG2h+OUgSgEZ6eZGTMhLauJ
dB3B210CqFvHRP1OuM4/HJehQZALp06AeUA6RqhKVEM/M6DOvBN9dlbdgBEv6H2WHgIL7DrV3u4N
u8e41Y7r03c0hvPa06fHzrHpiu3Fp6gjqF2kbOx3p0uEu/GdKBemIbvB15edCBBmwy1GdjjmkMVM
dHFo3+425hNv/IbtBr3DHfnHv406MSqbvIxA0GGa79wgR5Exo1aesBSaBbvAGFCtlu3Dys36P77M
ERvqedoIzF4TAFVXoZwl1ISJJHoT9/8F1ttbCFsXjAh8G7SlI29zUfmjZ3N7sUBLYpKaDjKZNi6n
T0gIKDIge2jYXPu/BmlatjH0MqsCci/IJjl/rZsnHiDqR3qo9YI8vN/eap9UF4gJVSZb7xslj9Bq
WAw47kVv0rwF0a1WWmSkyhaNxB3vIEh5PwBGlVzq4CLeFpdsdbUw61KVahbzbIju6sm6rT9WyOah
KDoIRzt1TaPazyUGRtw2v/FEJJIm5CXgHn5lvhLtIqA+O2hul/L+X5JOY6IKJq2iljU7950//xGu
4vObSTJtQMf712tEgUP3d1lVOO14sty1X83CaEEHIUAZjbHWK8VJ7OYVszLv/BVYxT9onrRpwSFR
5N47Nd4wNqGG8bQj2w5nMzzbtWijjw2RMJ4Su/zRgeMtH0DIpPGBSjra1ICP5DP/xjqIshdNLaIC
i314gUIA431S51I+xqJyzos3IaTF4g2pxWN1AlVJD+Rb+aW82hCB0CG3e4jOXq6hVYnKrs8+jsJ6
8nrwDBkvufHVNCIonrGBb3E4/g3gzC8s8gamUDYv3RFRP3jlyr0R6ajeWsHejsZ+Wj5xVp0Is7or
Dg+7dBQ/1Kgl5wc5C3sCTDPI+/xToMFNU/beJffdWsdnK/pWYCLTOqxKAjOzAZVwnLH7WRjKxPOb
aGp5+9FNqCARacDEZlYRozC+j8Y9oPUnZY/Vwu9DsE0+0n0uSufy5I2J+G4B1JQGoZ4lHiOrq3df
uO8VoX2Ma6pbrIncyM+Q/8LYh8QeqzYwmdZXkjpMYhPajUjdLZ3BXx4WWUliHRCWMIfggAv2Rc+b
PCnyftd7dljDKOSpeL09D/N/SYsKhieuy/i/qVrI9wAaBEF2L/eCh5E+xPTKIEN/ZtfRm41eX6K7
4VLEm/53H9U/r5cac1jr1aibC/YHYypVptonlrzI1cS9SItlkbOLxohYWV6mTo41bGrG0bTxZ6L9
gaxX2wvS0hgaToE+AJcGUP7CwoyedcBpykscd+4tkZA/apE56Mx7aaywv/H73EKyW2UDcOndp2Hs
WZBf1G2fD7UzBjU15cz+pd3E9sMH5JMOz6bTWlMhJzBk7XeP+4SZigaycyumNYnUdKYy1fa1rKbr
4Mbm6DU1tE38GDRHFoySA8MuHO8V65MLyvk23JTn8Ky2v1YRi35A6y3FY+y+8TCllLX6OoWLZJSA
dlUPsv8SfkiwMZuXAwpHrRuiYJg5hxiEdNnjkuKs/Ns2Ok63iCyU/04znZcxsfE14fx27aYdGy/+
YHCfO7v4WPJhuNdSsevhpdFsuFiicMPm4VWoaSGwU628t0YqZeTj62BKhWStOOKyELL3eJ5/EDL8
yUCY3hHYLjVbEVo/A0XTAXDyhNbL14+SlQ/sANvmHgF0PG2wFH3IHS5w+GnMvHjFbEqdsBGOInaj
niqoDtEgSaVhb7okCHYJcIKPHq7hNIwr4uQjsD2RZ5uJrqiGQJn6nVRVldiYToRBr3BAJGjmpIY0
nFRasDUBvFYQVnceH0EeMuekuzSZx0Hglq3nKSxQZOAKJhJnT/xA+NYCWtGWdIY3jyLOmHe5o51X
6xp/78xGXhVI7rcux2hzDu8q6dqN44GQ2k/zJcteRfrVeYSmyuafJPbaQdTeDto+oEsNzEjkb48u
ETInhhGU6Y0EJ/ErNhNe1/99KOIpC9Mmx7skla3c1lxdYKGCHpMIVmVibz63khtp4oBmD/sshRXu
HPgXC6leZb83g9n/HVoVxYsg/dhLZjVVp74dwuspm8MtT7ZjugLjKYFo9Iw0ITJ6lFM4j2h19wlx
JZXjy4m4k415pdF8Nt7uDOFEl6iS94fn7WQbVzzfEtRgkoYdhQ/AVr3YRVWtF06PqUOQwCp6Jg3+
RN55sOj35BxnKYRvGxX1DuO2u7stIYOirNUN/ic8TwikeCAUSZBIBg6Y/dozKm/KhIIGlGbj1L79
bdyiEd9jGJaSVNk0EidQNj+ZxW2inTgPI3YxSCMJRQF5LocRqMxSwZWkl8p88QDVBqQzgjOe5l2U
ln4XWnz4kUuw+MSX/5fOwuEFceqK9CqjZJh3sbliwXZIOmMIOq67kCZ142RjZzE80hz5eoY5gibP
9NB1I3nmO7ukXM5LOagdJwLrFJvwWQU3FB6PLe45QtJWbv7XtAqr1/Jel/dyizJpw4f1eM5wCokV
X0UMOFS+h3mHll1xGvudm8Hsu6JK3IF/7nyJnyDCw2GinefcqynxdWozGwHojMO9XLucavb2fJT4
nblSBfrloAKCm5hab2pwW6YuuYYC2bx79rzX96doX5ymwGhZWjY914oP6C8JllikPYfTP5586a5H
jdtkKsY2J48I0qlyMg5A41+64UubigzC5Fz+4bt6xSFK41uq7mKl8aQk5nUQydaT2lJsSNjfb1o/
3rV0utkT+8Z5REYSP2TpltLT6tc+jI1QQwWrez4Fwh2wRIj8GmPKgs+KSXaqVCjb2kg+IkhYUndi
v1M10XUB3VXTblWGMJWrbOm4GjdhE/JA9f2YFYv9CO0k9banGx51E4oJGACJu9cN7KyunWBlqma6
pDm7MwAAeLV4CXWL8O3/hU/QClDuiCpGBDiwbwlQJObkbrptT562YeXYQU7MIHqq7rW1nVGq2pBZ
Cnc4JUp8Q40TcZXQ/KthTWsGT0hoRxSdjGBfbLjRT1FW5ydXdE+6IiWMnL9APEk5gcvOO5AolyMy
tm2EXqaaDmDM+TvL6CsqGmtVYm1Hv4G1ApAWc2I6qjgnadBKDQFHSiwIBpctB5s34oZ2/iHp0PT4
BPa9PnDo31AQRfSLr/gPX2GazH3NCao4P/suTplY4qRnHTOw/M8j7rzUh7XyK94mdO2MxJKqIWEW
XgXO0PL+M8bnyEr/ZtPQy7BMYkY66QUsA1nRgi0lVlw31wtrGqSCXRYAdxTAQFPVoCXUTNt8x4YT
A6igWC+HJCSwWGAvbHRIWTw++R1Hb/8mtfVlSW5vcMXSdfNjypwmuiETaZIrRVIncaja+0Gemn/n
ZLKq1uFDxKiVap9qbfJTP5Zqg5tONIGncKQl9pa33uxkx9mSuGt69GNuXp6rWvBOG8goxDV+5Uzf
p6mXkwRYVyckmCloBZKmykaSw089u0UmK8Va1Vi1wAo5PGUWqk4sOLNtlqkaNJ6t1PrPSFgPaiNM
vq4wjdDMhJFhp7jHnYiiquwckHsCgHp3yAM5m6AKpcFHKSb5oX250uxOY2eIYfe2WUtEC44rpOK5
ZErha+3BhZPgnkh8sTx8vCxvw/oe2ooH3ZJDpSETx+4K6zekHn40XD8Vq+37I3yqs4puwlA0jZBF
OtiK/dxZOuBk5SgF9NwsEnVwdZdKeVbQA447RcnXSXJBP1DgdgUddWpJ6JlA2YYoT25zq6NvKLsw
G8gE5fJRhjNa9tfWlFu+Kd0uFAeU2kjP/aqSJVBWf/Jvn7ov1/iyu7X1ys9x6aj1bFeKD3PouA4i
zMqCZkksy0q1+ZZQEJbl5zQ/AkJdg6tyiDSjvejK5Q90us8VePXAfKfGQI9LUTM91XiHlvLftghc
2zio34QIamKzmPca0wfphhKy0QyYw1xJGe3bTrwviIUJPsosq/WIg1mLtLqF5Xnu966mONwB6MDI
zMD3aCPJ5ZJC+54aLVX6aThA5gsWdHVOV1/8xzPuZNfZkTO0MpcMBQ/kblVBE55A0d2S6LzqS6ji
cg0EYPYJlMN5Air1f20KXaKcB76EcSPn4DGMEKTicIvdvlVef86aV+hcoeWfGvaRQUvTovItkXMb
WrhIy8jb+t+gLSi4bHj2bbuYb+mD7tm0j99ITEKGEn0VkjyZJeevU49pMO9uNDwCe5NgTMxBrWkO
UGlrvVTVP2h1wGnKJfq6ffWQprN9hYF/AUzsDdw3TqcUcguUcd/Z/3lfdNtu/mzwuzvTcmL+xck9
jPXiOCgCNeCpHwMez15UIb5v4ldyii02wmvjVKG87u1mM+hLs04yVXVPwodgrRkODlWOvOLQyYQB
KqX+uOX47Oe3T3sTKePM8PrXllWZCiqmSJtU/QoItWNEZXoBLO27ZT+xtKsZzZTHxvejif/JS3pA
M84oucXXOkBi1SEchgwNOSmbf7bsvdyWrOqZhMokEgEtNc37mfuMBTC7r+QJt5yqr2+kid2G5Hr+
TSxk6Y54pQ0jqr57qaCCRxlSv5fUN6i0iDQilJ/cPXxLBvFwMjFbhkGIKgKlPQlJ4MZgV0uJyxtx
D3sgySDT+tGRWCfsllP19gw9lO8TmkHcup8jYeFS5YPBq/IjAXwcLeOJkpkcY/iRP9dPjlZnmCm5
h005rudhStePszY5IT4GiG0tIC+Ua1GSr8ORkCAmFX0zHyA4cVYnvMzNYLvIKyvh7HLdcjgkjylG
0j8JyK309vcEZoIiMl9Rc4K8EG1FptGKb3mSazU9NjlxL+12h0P1MW2dUODgpAKsFyMopEhZFxRM
yrVwmCMDexxlMp3l/gwMVsW7D3LgG1ck25cS6p3//vovqr+zbLMt7qf40Wh5FjiF0vUVL47Psnrx
F4JTaM1AMzJb5wPPDmP2NGwROlu9dzD+fUxMCmvWT0PeUPZB/W89pdZGbVQ4dtp3OCMerx5Vvg/I
aB0E37eSRwBrZ1BwcqYoKdTehHolSpi97RTKb3dfMqSAjNmsYouyBc+mCDXBIYrvwClR5oX+kd7k
tD2fBccmy3S9J2nF9aOvqX3C2jNQzT50S9jaaCUEh7U4hgfGq0uZlOJDLW8GcMDTyq3cslecElLB
F7DyUtTv/SmtmOpMoXa/+EZUlh+R/u3AXYH6TkjFB/IXd6AM1Dl8NHBGWyBgd9FwkzWWC3c0/jWM
AFaOzErXfnNMYxY5qBZHS1+gH8e9CcBABgBjVbKLnuctxPS8bWNm/FBN/4aXfKNMQcA+S0M9zjkM
TJuLy26bNCa1w2XTWht67BRWFhJmvde7mP1a+jqYH5ZietDdygvRy5gB0CzsgC3nvaPCswvsNVlf
nMreu+vaLPbMr8QgwIhhNN6zxM6huWPwmuf7zAZyTMpUzLrfCY4WEGWQYM3sY00LrQd89vl/AhBe
ZQLYRM2EfsZoqlm22soGSnYKXi505/n6Xk8lS9QsYC+5+6IQSJlGAdpUKTgXtbJ/9ie69y4y2Nac
4iEcGf9vb3HDGBU9KhOITgG/Ht6KuXpVZy7/qaT8zvMMeeBkTdEvrQaB20wryEySuPGdXWz/iJ0g
OU5QlGNekCyG2lDvYSm5m0UoxD/8QBzTRP1YWqw7ojlRE8m2lvgSet+0oQzKRiRE/Gqb/LrkPCpa
yfu+041KJAzDy0F5uy0M/5Pf8nMz2LoJiOdXdqYwtdcPROcLKACcUkVgnVoHdDgDwzem6jsS/2RG
RGN8W4c+Y+KXXgIJPrbmX2SInXoaJX8AOJsf1O5nYA+2Pe7HNAo/he7KtYBkthWed/WU6Md2O6uF
Uk1jLHO7t5zdDN5xZTNdQXdMXvNdpUqIytzABNYVvgq2jrDMjRwZymm9PqAc+3jYBeDNoKNkSwhL
KMRgbXHaRK/2S1bWrwKArQZSGgUyduT1SwQAACOPBtETYZXqa+od4P8jZwaX1YUJIDbB+up4H3z7
S+udGE+RN8UIROf82c89whEqcpdZOiYA8GgtnbfaVvATXOCOjJzhHpqklSo3pOZctYVC0rJ8TBAU
syQLQNnJH2nqGuyz7UUpv4MFRzPij4z3S1CI9OhYMpjLDk6nex8OB29LtDFnDS6XNf22TSSb72yt
2qV/pjt3htXe239//aH/B76Fl2EQ2GxgcpV36YAnz/Qrnql74oU+s76c4pa+5/vUJDPao4N6C+zJ
UAvf5CrqAI8fWcZfMhQfNuaoZwYblhIxMpBHo21/7UgD+E9TKT5L9r1Hy5FiGNFVcMZdrFymdF5Q
AGXvb1fl3/uAVTaUcRy+6h7zarN8yTIOW+2TtUB+gD9nS2T0kTrYVJNu68uGee33hUge8eqUvVkY
nSV/XtuVlsDDGc7KDRn4npRQMWTWarP8dNbHumHBdbuDZWLqfOl+ttgYq78SvHEhWT1y5AGe672L
WiSiKgEsYLt02cWnfu1PDSL/z2qjL9FJeexZ1/p/qCeATSfgbePK8bj4lz5DRHV2R6MOBaDpp6wY
UhJSefvPMRkEIDJC0x0QYt23Zrsprbo1JeHPpQY3/OIitj0jpX7JnKB3SHHNcWB+FzU8rCtettYs
FPtMyEAAyPLQNiz42FXuwa++gEPQij9H1NTx6sZ7e8gpnhTyS76uAP265wIej+xvpeKlhK1VtNkG
XXGooQWw2retGNEEbBpf+jGGSYBTaLwltgS4eRq1U7pdxJYYZ1Qo937/Wbx+x5PP2auYTAGT9xAL
8bXshaq1y98HE7JIx/ANiTPO2q3hZYphIe+JhqFjzyt4r7m8Tbh6tmxwQ6fFS5Iooss5kLrjK8m4
eoqPvbSfomB5Pv8webQrqq8MbA1fLqaMCOYfijYrJZLUOlduHbCfM85f6ap3C2LlWbXtGnXOQbgd
tMv09Mw09wt38VnIrUYDo9WeEzp7Yik28DSP840S3YEAfZoUPkOWZNz1CBSGYCe400KGest5k8EA
NNKBqYCICe33NShPe/pqBpjWIM5b8LOjPwnyFHmhkDi8n35en/tckFeD/I/TNTfZtCzOA7rW5SP+
2GdisdVBlU7QhosHvHvGAJv11JUrB6b6g8NrLOAQRN+raBl4sVZZx3Y3eY0vijo7X3WQNqDyRNdU
/XXXTy21JVjHmcSFaAG8vGkFqcGOnaSxJ1McnzGMoQuCx0nZjJipRs86IDwAc2J9+y/5i4pENib3
QbYFkAuDhk1awonkV2Vmi2xTkmUL522reUNK76sVsLlzA0G/gyA/aGJmV6MFROqaAdG1E8Zz/3l4
2HIiIws7gOVwjBZiOKSWSlvIMT6aMEr2W+e6DiYUwkphFXot0I1nBl+h34k0KEHG1JF0V/CmJ0W8
w79dk1KyjckBLkz8BDUneiarWCJaCGTjeQ0dg3TpQjtNCVMcinWmq0llVSH+TRC7cuViHfBCciug
GO7vt8GyLDV7AvhycjXtjus83Abskl4q4YsrtvCw+2+YFxFUdHbW8QOteF6zF2LgHEos69yUweep
brGQzYb5MeXF19J0jJgB+9/t7w82ktMd9+OamU1wBAC3GXtatg6VgLRL7pi4Np4rfJoUMBjoM13L
mIE54YpqeThaHDXbE/kXJ+U6XY3EYFpVm+twNmVn7D/FTQDiqaPJSEpHzGFTnL3xMwpY81Q3vDr+
CqGIXlbduO3l5OSe5CN9LjgcLlTa8X6LwyHeSHAAcC7HhjQrrZ/hv6yHULKh95utsFikNd3QLeZw
A/e/SWDU7Wg3rzAIaJJGDlV0YMS0syga8cjxb750eu790Ur0Asu7xFH4IU6Tf0U+zQTwe+/O/5Xu
7o7q9NAx7cAPduyFYtlT0ZVqmwZZRbpTdevNEMILtTmlODJYJBXloXGawaTatZpszqQNvxfeQfBy
+qoj3uCfmwbNiUAk/0hFnOS7nT5vZ38U5NRnsUaICYvNsw0IMyNX5fsUhapULYApBmkq8Me8lULX
Zazw1XhaACSWJPgtlMIJNT0iXMjgXC6/4LP/sF9vQizO/xmiWOk3QAQdcAjJ1MKUQNJP6mM2XACU
cebHlpynQqdOw7qsST7Gthwwd7hSs0dvUamMsOuMKoSyXMLsbnBbeUheK2U6/eZ8LyUWh2M0lJNF
hx6C1YQBnDd3SwCKQ9IJjms+boIZwi3CiBZk+NzYmlld/Oriwsum1P4hur0FUSjEo0FQ2FlW1oQG
nTMbnb/3mMzFun5fj2YHxsgKiUyvIXpkcIvSmQOaLYwm9gm0Q+ZQXdZ4zoouBRYRZTAsBzPeJtTH
vlcJv9kHXxj9Lm0K0Nwo5r7VAh4nLRf1fYKRQa3GvFcPCt6P4funsFc5IuaEiT+XPBPUUOdQfVf7
uH5IlQokUIrBVBO+H8OXHS++M75W+/I1NHHUaQeU5u/4YQ15q+MYxHZrQjI0x2Sl6cvFIGI2g0ks
ArxMyruVu+WY7zqeJ7vbqU3lyn1yrr1EVwEYMHDBq1o3sJgrowjJe06aMyd2lDJ6ieS1rvmNH7UW
5WwHOtuLyZJGkaVzSbHeLQJzYBwDDcH8wJ4fzS93VL6eWdH5rySPRZ+uEAmRHVfC/o4PqMWcfMIi
wv/pfOPYg708clgTfTxy2KWU0YPU/0LTe3nG+OFa232nx9oTXZmHAFjsoYAHB4du85xLfURz3ysd
7CkvSIS1Kv+29saxzGXe585w9h+wn3E5x4w0pxTmaTPFMh9PgeBjLs3lGDPy1h29Xo4el2ZCIkqf
IXIHg/EcElKUgGC5dnEQFl6AMqE0c7aTrBlg74MtEnIZSw6ZliEhndJCb1bkpIH5RlrWHZKhAiDo
pdFx4dJ9VN8LN79XmRBVKMODmzF61YIP+KJJwAKuWDJXjeJ7LQ6U7zZfmc1ocY9IX7PsOTMfLwJv
FmqD3KXJQ5XwzrsEDJ6+1ozdOBKy5KPYckpNsU2JOePRQ52kHZ/ijQs5PiOUQZslI5gS8CaUVCzA
3KcHGE5fOTIDA0VXABDU4L9vS/IC/2X74650VISpWx+k6DZLSm+OAmoskaXraKJaKyFIV5lOWT37
bdt+iL3KXkqcbzAvz/Vd5mVyDdUJBP/vEb/pXP0Z/i1Px9X14cMpCpM+pYoeLszRi8s3vBU9moF1
dYaV1c4YGz0+/Q53WwVoc8Cb+FlAcbuheaeFPTVKyf051pgoH6tnJgnKdsNjmgHZTYYHPvIeWK4T
tUqlpYvmy7zm7m19iznB8OW4BSYWr8IoB8Z6XKYJHkSt+qDkw8r4waMFxJ0keauPfc/fgt7rVep+
hH7y44YS9L2I3C2ifvBW8MXetnLeszQgJIBp9JZJzMJFv5gNWu3ZmbjacyiZ+NWwehw8++GiGJVf
yt5IzVVGvUUXqQ9ABZAjkNuqkITtq17EcmjYr4uaPvBtN3AN0N4/+fCKeMGg9USP40j2lDt2UicD
WXgoNfXwkzptighxt3BF/d/QKST1BXxa4+nUmhWmG/LUbom3McvjN7OZZMA2HGiW37CsrGOPKPiS
6gV4qnK4O0ZKC9ekipbMr3x0QFeYz0j6UYZZW3k9BPPAeabKSq9SybEeyvP7vSaf+Tdb4VX/zGQD
BFkTCMzBevWc3H81URIqyykiNCVIfx/oficjHClgUaoZkw0OlkpLxf4Rv4ylJpUaXQKHH2mAFGmD
qstDfL1Ue7S4PnaVSfAkSLhhBwqU+Bk1bxMG9XdjhGEF2ytZsO3K99G5kVhqJHocuZBXGuMx3q3r
anCmf6Ay/K35vFeEC/qkQNWEjI6ydb/fZXh3NVshOHhTM9ntetnE1fSotPqsz0V/l3sZ6WqeesSB
YatD5S1gLaXUOv1uBoijpvJD1pvDEWN8FU7iNrJ8Hi8btSEn45NhH3aTj5B7Jo3H6XLzy/FUIST0
ZhzOehDfgJpEI++/+CuDa/rwUWPQVSSK+k8vihndgD2RrwpPPfKnWDxrZEo+Po7MBgstIbAvN2On
Qd71TTZ6ipyIHbYvKUKlYUUJBqZb4kJvyu6vT/Z0UbBgwurTOTDdA/rxuW6DpGRg3NaZpxO6/zCE
ts06zb4aqOHhu/ijiHGWYxSSkJMFJ2of+x8o1t0JVAR2o+zciJ2L2TnuVY/HekCM3Y0jjUBB+94f
1JeV/2IkTUWhlOMq76SzCOhMKA0f5bK7tcDkPrdn7WoFN4gU48nse8XlO+r33RddgN57NbfEnPaI
pIYz9n5qhBMEiYdvM4wH1B6QaLCK85UmqlQEFbd5Rd5cpx5NIP4GOAx9lVaB3Ury8ndxlP77DqAT
HJ4SNlpOLCdWWBD5APHMgKAz0bx4+t54DcLVtgSWQgFRkq5zHuLmAftExCcL/Z6naZ4peFO2V7zl
Uo/wqUqY3MorQbi/wVSpGcb1EKZsmohBgg8p64VzozrCeeV77fyiGXqLn0viIHsxyGCboPjv+dK6
JwTZgetjy8dmp8VGQniSyVnAfXAoHDVonmS1SvmNYa469DwASjl7DRSbVMzOqOLYpV+242N/FyKz
sU+kr3HHludXLt/BjUixDCwg3AQj0Grm/lwr+2KFT4WPKczbYVjupaKl5IsQM5Z92sFFFfDLXNlW
UVFhMlD9l5wfVcIxOALb+GwUainzFVYW41puTcx+wUZeUHeHOQJG79Ke977BU6vD/zC95z7AptSl
MHXOGpvRNmZf4Yoov6a+Ln6POgXt9nbc/OnTtJIt+2rozfeAqlbU48x1KFkYPzLx5Qj/5pIHRDTk
U8rxCLkyPOWHQZFn2W1EXIN9gLQP2KNreXZNE6OCsn5ZiVVOSPGs0bSPBbp0cAqovAC1f4b9qkIh
AShhWzbjlr7pTSz6eSpY0U+UORzGKoOgiYXfsuUwr63RVM9gf1Rj4PUoaXHGEXF+2ZR1/sGQspd6
PR5cVGBunIn/Koruwm/WmBiH6smjS2nJfDRKuEKaucIABHV+baQLrIYva7cTtqeo2oG1ESFwGW46
TqVPPQLFJgmWLDuBU2LKtqijDAbGHc//2ck+aPB0UVtLVKrl6yOsuMN67nUakW1WmikRQFfOfjIa
HxrIaisL2WOlPJgWO02i2HjvfsXJ0xZUa/UqYgYMoZqUUqUnzH8mUEv96QrpXOck9Z90fAGr5hjk
yNqApbmWTgsTSmtPtd7NXj1BJ79UTsozJqVuq4fyyUHs7Bf4EXSVdqSUKDWTx/IedrmHwq3OuZoY
UAq/egrRzCyQc3kJU77sXGeeDJVgvVPlpVs6i+i6NRN/0N3znqWBWuorsEHph06qa5icKalIIA8k
L3hjXxjf3GQftx5yevvAHzg6BYDuiSppgqMC1jjzTh15HvZ2Zb3UHiKtcyH8xHOu+erNH+lFhuD/
fEEkkHEz6NtBYXSU6nBxOkcmFVZCyWHy0RAlxZ+NmMALg4RTTijxoHIW57VOm38zk1pmazmkSn50
fqn2YbqyQqqfbZckQI0lcGEit1RauYGGbRoYxivrvhMdwuR8QevFm2tdoVCQYQ4ReZwgSz7+I7Dl
/IfcAdJIibnS4XjjlyAqMOSc5ws4aCuf05sogh6LJQbA+rnXcvwfp7jsRXV7FqVjJWcFV4XQEwf6
/2FrJag/6Sp7iYeCzafrbuMADyLHTFxyQPjlLYf2Tsu4hpvQ9Rl6KBZ32Ao55hzGGV6CAgAgEyCg
0NgGx3TMdUhF6XFX086/Ywp9sFB15D5EoH+n15EXYgB4vaf1BITSx0KAyKlXqCiESox0VD6tUzBO
kcl2DFKz5uJlN1lUbmdfuarpsqVQ2Xb4JizfirUH1r9PVgBZv1gsHW43XGm3Bi3m2+ltSpFt0IyC
xIH9Muy25hvg8UE3fktodhwZQIKGIxzomDIn+UR88U6TR8h0/crObzBZbKeBXoj3+01Z6lAsVTfW
ZNV850NS59zEcs8tFD8h2NaAmd4mEbqt3NdcXTnzYoU5iRoVzbyjRQO2XiUdNmLMoxK8RkgrQJty
abo3nGATkGb2AOxGyqj2RECW1PoWjQ9HET51WiMRHR0u/BHbR50QZIEkVyThwTlERqIviZ7Nf7uD
8N1einfyMKC4Jje46C2ogSyRQK9eirtviyjdk3RSl+AceS6sq0AFHzmLoBoF8fOgbdiy05yYNpNN
sAiTNJdYl6A8GUFEAmAejJ2+tgyvPvYHqGBS1+WWpdDI9yPggspH6UpD8z+iIG6LR4dkrxWWev0+
RyWtBGrOfoo1fsSxFFJ/KhyYYF8XIvYRBrzsQRUiSQZHBv+G34QdxnR5ZWCzIDdb8sdxWZh2PJIb
IDTBh1MYZradJvRspA9mZ6F1aMk2/4CebeNAl5g9f7b5fYKCoA0rCCqNuDI1YCjYn+rSZkrBsNB3
+OPOmoxlLBGdYnvzHxKlCWLmLbrsFJTvZh898vYzLUkMa3oL2Um5bZx1x2qeVpzL2Jux+H26lMdi
INAdnukmsjB2Jfnyr3kTyWmgnVeozqHxG7Zy9acNfn6birgNUwLk1vbU+fEhtuhokxiSGrzGxgcD
8F6HkHZ1IwuOBH7W7kaTZ/HDq0MhfKSbvxdet3XYVrO+kx/uQ+3od9e1TDgVb1UVbnJYqtYbgY2J
VlzneYHqYqS4mj25JojIJ9AATgYsZ7vCLxDHe7gbhyQgLdunMvVpwfmUL49tST4cHh/U0T2gRQBB
zg7wL/EY1Hgj3lUWy/oJG2GhTH+snw6ZtxTCV4vYaBFuvAeYuWGR21QleX79K31LBtpYIH9Hou50
zqa/8JIVejWORvAPmuxGgJb0GbHe9JfUlmT3HU2sEKrHSQPl1aS5+rbE9L9o2C9uPE1DNVDHziQM
asoleHq18aYZL2WldHmaKKSAbsil0xwsp2obABmSsPuYYCl67dOu2BKgGQ941qoiR6ZM4qVDGUhB
jP+7ftlyai28BEsu/RPK/ZSKTQkuWmlCpN1e/VpHwiBL4mZ9HN9BN7mnCPjtKwtfJk6LrD2mQQU/
gArZvYnt0FBCG8BW0cqM+n1pffe+GQbZvgDgXB2b5K+RNUbgP21DktMuwKwjdN6MWwfrERfJM9h6
R1iofGI19f0e3S0MVtM/eTGy/zjgRo0JpmVbpYf2azhmmQtm56mjPqOGUUKK1AxsXFhJDAv0O2oi
+ih58cS1dfOCHOvWMemWLe19lvCjPfBCCf1yUnm/o5FY3LhDdmGMdB6Zg8Gd96dvtGy2HE6xm6Pt
ZGQFxa9u4ZvcTQCXAwPl+/d9grGcA07WGjNfGCltuY9bh0sqwIevG/ixUBKweCAJJZz9GYkMTWfX
Twl/6ICfAfcCKzhl7fyO6nXYt1Ef0EM2NemNTy37nzsNeGS7WntBEOBmnwtbiydJEee/WBPAGbG0
pKP5BGooMibLTi4DVrtH2ayHADqUDwKKgoc4Zii2pjjIQ7ByJYDSNCwKrgKHe1lJCqNxPg7FOjvY
7FWXAVQiQTEDEvCoU4Arl1SHWCarE39A3dA5tQprb1FDMExEt42goIDQxatRClc24rm99XPMW/w9
cteO7vB+3vOqYdwh361EO2YGw2WhV/h1FhARAl1zD39r2g0EGnwS2ej3N1Rgt3UhijgrUwb0iG0/
pukzb9fChf5Y72UWbnWSrPSH2e6LibS1dnJrxUfIcARnVz9k5dAoOAZz8+wXpl1B9FrSNn4/FdHH
orlyEiHz3RKL++8L6vBmZ7gL2FSD/3ote4WC5zP/nRnAc1kb6FajMSDJgFA44aZ9M+/8fp4QkInT
v0dkilbPcgu8i5CI/Janov3/v934kZ4rs75RbsI4A2N4iV2lvaTRuc9FyuY1TGsM5FwTGrlGry6Z
0y3oemBItGOKB4flXcnuSTCijnLf1nDgMmIRfqtk6FrUWfFdRgI4bnB6r5HLPFPld/3dydRuynZR
P1qi8swNbhv2ngy2Zol1eKRWSL/t4HXKrwt5d3K26MWa18nY24xz60KSgJ3Su1CUFB3wIxBRRqi/
KelTn3MgEDBt6bfxioEbWyz5fNfqR/ZJ6+lIj+we+kznk572AG2F5NwDPyjVdbVtxHP04m5Pe9oF
nm6mmQ+l8BXyYvSvHeVOa0NfKuUIAHiVxT8ncZVxVOUEpMQTtl/PoxnTdnOULsAMETIZ5gU8Odq3
roKG2LG0EDkA4PzMDeyk8QSuM2ZNIgEq9XHyh8CKMByGPPwlHrIJgb0fePcfQHs3q+rZvvJXCfgq
5G/KXUCCTyxrRpbIVVv5nKGhGnVTURB/vFbjWksLHCzDE/TQzCgTkGuBJfi7C3RwYVBznPZxFLbm
RNeOVRfF4rEPldu8ULU2shuZzYFh+bm9IcuLAysv3X1V+Ivv/jxovlIf7dKA2igOwfAnyBdb8N8m
kZzZ26s35QuFggNilJzx4SiKrCDDMMme0XKAjfCtoUAAhbn6mzPG6OBe41DVyex8rCs00aQL+qmR
e+uinFpb4lHX6Ls3mG+BepR6hE+1IJphyokATxWkg7c0Cnx3hCaTNTLsxRPVCLKhbWqAukEvSVgg
YvwklPuJJZU3cruaV57Oa6f8dPTNafDrsr3Ve06pPeifE2ZxBojEB1VrJMT8OaMlGsINW1el6B4b
mkRJ4ebO6yB2jaWoSogvgxY+mZujT9FcNhWdovgRISzoQGJmvkYmZDSoVrpDlFLD3qNrnPgecMPT
31MWRTwVur747xaIg+euvFj+B1lj8um6AVVqYbDRu8SNM/lCGO28rwJL7291FVbyFNP/b4/oiZxd
bbF0gjKkbOXmSdEaR71koYwKUJ9Y51IexLdR+tlmy3GM+m8/yXmVSXvK0WrvpOD+eAwacan61LgK
OklhOTIyffFsKH1eDoUr0myuRJnHCmJbSnqzHutDicM/SqQXn47qfNHrO0xgifg8Qnxjmoiwfglq
ZsevbNBq7K+9DoIUXGItta8XcZVJX6W3S4apbcx55h6S9BT6Bqjh4yZi2d61h9ly+Egv/nkSyey6
WAiEDLDVIeTFNejeGWvQGWoL8LsLmlzN8s6xO3Z+ikdLeEWj13njjh7gngUIpeU18MgKmCE9J9J4
nPdtdxjgT6JJk1HL7q2Ga5pq4nOxInCQJnjF3K6vzNoyNGqaDGWn7g+UBK1Q5vDi6zWaD7dIVu5r
QYCjdRzKf6Y8rq0ZEABcvHD+JqcrAvGMyDlToCgBa0hyvhC3R+QBapVO8Urg+hbprTD9N0K0kM4J
Tq8be3pttC8imu1n2uQ9OaPHpvakZIuKJUGSi+rRkCx/k9oaGC0Eb9G1WMW3RMOTU7oz1rVY/wah
kuncec3oYbLdWAFS6NLZXrNQXwKS0G8UoRONUqFOVwowsrxSOJBcxRSAys7yxyc4OTjriqKHcGAq
Ajnu3y7fzNHTosRnBweEfLvJFNzDEhRc83mjRwNxA1mbPkZIentpceGVXKeDS45Ijq7tsF+x+Awk
vryckips0HLYB4UuMQr/pXGtC9pu0EwOHlckQqCp8+5j44oXKfKpCye7BSgTOgi5dcfmIBmq+Nac
pUSbTos5ghemClUuwSNQ4fHzQi07x8ukH37YxImKWCGqicUXnY7XzwtZRWSb5ky1ZlgKWsSxdH65
Udksa/eYL9Kkiv1wgrPkJbujdHs0o1c81it9Aaw1epGMmTUha2WHAX3p7KReJgZZbQf/DTUAmXVN
08RnXY+LEEiKg2XHiu/3N6I2BGWxQKmVfGoh05mmV1ugoP68xbMsEnjbXUS0UY+om/nqUmggU78D
rPYm9dVAbQy/izDeWJDJM9tqRCF1MY7CnmKkTfgevZnXsFmwksyUvIdr32W1XUBmWBG33gTZDEzR
+duKOMCU99wMigeGSOpeCmJdXuId6gfYEN7SAbIhCw2rSQ/DvylqAyMmgxsdXtxFQTtAsdLS4zHz
YL4tBnHjJ3qwYNHL1FfWb4r/kPGOxvnQHj4BC//r3aXPllZ71FkKnOUeaao2sBo+QzrWsOecoyaX
GKL1id5BFHc+WTkhMT9NwouSwjSXhoHABZnLV1AZe+HW2MgZG+wGBkHLwKzaU7vbSX6xERVmjVWG
QrcWgKN20VC5C48qj3O9kVCEKdfOEphdMbMv2BeW3xI6p6pq+IE0AdgjPeFMteLgtIYdWJmyX8xX
06sVzOMmQNVYrjb2TWZ+XvX5OqoIrhJycQZr+KZrKrXdLn1okMx/xcVGPRFIumsZtkL6Zpr+Y3Or
6GO/UhwajbZaei05OkmJCRe/MT0b5+DGKoz100n2Y+xIsNVPAovTV+TC9MlRGdT2jtG/IG3Di/Ro
jKac41gyaFBDF0Nm9pAKjw2vIGO/NYdRQiee4PLkXa9C16NM6G5XoIGPugYNVEr/3TxFhY5A84tN
/w1Gdi1OlVdNUrIcQ74BHbwDbqEhqmJuR8QXmjU4H92syc+nrzeJ+8cWYBew21aEw2Ii89Dfh+sH
70mXKFFvcwWdccOws9DE9mJTDkRhpykBPFKGb+vJNIDKiU2HkM/zf4OPxydG+QziO1mOrQBqwc+M
8UGiXWkK82Judp4rPLcPM4g7u76bsMFVw+qA95xj4ukzY3gmZwLbFV5UXbxAHw0cRlQVp6vJSYGF
UnLsIkEsD2P8CwcUWkB5BhWmCek58Lrdpfk2ox44L20jRB+G3WvHScoDfP6wArl8fMOU8Viu9JDz
ShUMvwFrJJsuj/hK9IXU47RNrjjXKeFr7zq7bHdkV07ssTtnf5aWNE0mUAXQpP7ypvRlLTMCwmGG
5c4diEfgQFZwXsdNWH+G5OnofZI+T6AV6SU3Jh1LLEqSlXC+h+6CWJYsE0qSnRAPtJqe5aVMpvDW
yKeka6q2JEqnQpqpCZZUoez4Bk1Dj0pWLyeuMNNXSkqAitDMXQ6MRr3QcqbSgUS1z7rpnZNcuJxJ
yXy7wBRYnsNlqwjEGnurWzMMFE80Ky17SCw7W7r+H6HiQA2CILEfdeUlX6bq3C23D8Twl9eJOt2E
GfZ39xzM5tSDih27env7wVq0aAXOmEsNt83kJTyXUvN6cey6e5OowdIdJ6gHkq7Eyy1MLw5/rJ1l
oX3K1kCZOw248YrwOxMd5eFgLwrW1keiaAuygaBZTqmVY3I+wd2rVnhCAhKTWWXaQ9OipU8fOHNd
8b9Z4JP4EcjdTP8BL5y8vIDb6jE6nt8QeMITNh4Jfn9p6BP/s7egjZGz4CnaxkA+DjZsuoguFakT
QL7wpKocb+6rdqgIGR+r7W5cZZrt38j9Csf6T4XDtX1V87ZwLLp/QAkzSRYr0zRVwrfBzyPIj/ef
79tDnHmSKffk4gegC60WGOP3MQLcV+ToRAiwz2gMiT3zwdV2jIAB6c6XcC7lhxcpX3kPjrGT0oTD
HcIXZZB62skrKmnX1hSRR+/1ZYDC4usB0ijHCbngiuot9k924F466OyAslw/+XZADk0U4GE8JXjV
za70vcpaLXyPE7bSleSRxSipXP63ADgYt8BcwXm7Wr8xZSoUPtqlZH5lDwW0znPRsnW4PcJ8ZiBi
NTIjun1JZY2C+dEK/itmLEEcTZZdz901M0dabsLDIX7FHI0dzjEEHPgD/dP4qk4HwpagER8+p+eY
53HR9cpm/tue98kfwymMqMYfkSCMuvICY9jUA2923i1B5+l4nb2lvaVepChaEm/ggAosJmWu5WiH
KOizwfDgKpww9zOdbgjRFc/dw5N2PJXj0Kd2l1gtTLydwyuQLFKeXmruB2L6SrNE/0mUK28pdLIP
0y1eGsQX+Cd2MK3B+/cVsExSOIas9JQxkM4gYp+HtC1P9tnwmTv84limc0eY3XGNo8wL5xBaBaDo
Uew4UkJUfyieh+RoCnyeBGMAJMzXlsUBWKi700Nb1C7PBwLNcfAN4UPBJnncD4XjzkbWtB0Jkm6P
2OdMdGFpPtSs2ZEQ9CPf7aKn/a3O+twY31EuXE18hk/oTGRXQK/hq52reejY0mw+KqmMrXEJVcMh
1FENKMWgG+OFTQFhTgfsDlXK9++R//vlpE1PLK94Z6apXiYtot21AsrIAQTXecxICQzaShLM4u+A
S9xptDpI98CBOcHId6fm2Fioa5YVUlkM4u/0jx8QT9SsvYzL1WLXnvrxReeVkVlb5tVlMOejkkK1
k8eatrXA8pGdBSNj1Yh86QE/J7qm36kGEXd5491rWrUOHoUtm3gFwDDlg4H8R0Gn9XwQr8NjnYP1
Kc8U6hSKAKOTqruGpePD4oYG9fagUn3X6wo0s4FIwfLu3lX608cAb4XzGpCGOhIj0NxOLGcbJHag
MlYKG3xsHNt3JCjnw9FEjrLHfiZV+Xvl7jIvUAhiSMsUsMHEDUFwFfxwwHVs5ikrdYLq/mop2Ywo
xkVUe9pGw2yUpNi/JAA1e/gPhaqDQ5OhVbPtAZgGgUG1JDi8FnaOdhqc4S7hri1ygXvpdGCQTFIu
LXvJMkJfzDMfc0FidYJ2/Bmhria705Av4+jVMKe4aYeqDPbUM6v6QPYvb+GXKbzQ8ctoQgi6l2SQ
/dbwWEp+FiHb7vW2B2q+7zLBnr39ekpL6i0PtX18XlR11T/ysFOfwyKqykDyXhN6REq1V5/oPRtv
j9kRMcYqutWI07soR8QAA9Q3+SfbOdkOC1Zefp4Ye6fhylXn0i4CIdGaYNvRvmJ/x9IJkLU4yKDL
bCgua4giX0I6ViBNX8rcQDK8Szd5Ik5geVveuMqfAEBUJ6jrBRe0ny+t8zXl6C6eVcWS3DKzDkxj
7zjTFRe2dt0OthN5QSlTAxqoyAEgA+pZGlGnOIJNsEi3z3lDdBQqrxOQ8fT7sMerpbgMrA5WHItf
7ctxTaR+tZWD3a/wLp5s7w3AuFDy2WVZSvpL9SwPga4kL9lWS8XgrsSzeDGiHI6A8pLjZ1aV/WUP
K9qc+LXsGPcoXSbneXvzWkXA+cIlPcysgPJdSxpJalLTCcPBRTcLGhvNPCd/F92vArdpHelICrCk
5KbjxsJvGsxHPCU2OMEgBw3bE7kUMycT2o21h0KdoksjOgXbhM+kIciHHngVZsa107wh7/nB0gti
SDT8WJ4YZG0kBO/sg/f3UCTC4cW3veR3tSJJ71XFIS/SIYZMs7UHDSrglMM0NNoLuxba93c9sodO
bca136fFJRxOrbNeBDUI4Hs3Ydr6tixkLxB81RZybcD7d/rmEmIVQQw6dySMBAteX0RRhGrDSHRL
CP1nkmwXk2JUsCIHErGtUuNZ+N9/WhVmHfLsK4qE69aoax1gE3sehy6ZG7uo1LDZUtUd7qce1sxo
K+UaG4p3UP3W3Gl+f/vJ3gjUFbnUUDj0TpLOzW8g2WKb6mgYrFEdPDIezuhlpm/Q7cYqPK2hcgHf
7hYflQMTZ37OsFSDWcpEXe4KzHoI3YTfUxiNXBCK+cc+o5gjLAK6b34QAMWjfw4gNMn4dS0ZtPuM
S2YJ20KSbAVxcVHKs6DrXjdunHbwO4sueAN51mwZuI8G+8x1RyHIrepOKxz/2D+jao670F6QbPx+
0wRGg7qTZY15SWXiuyQ4L1jgazV6gf/VgTAD5s9hUX9N3nC2/GrRwWSQKBn23SViGu6v2W32Sb6O
nIPXMRZ/hwlztXM2Ia2IOYeoTB+cJoLxDlN+Wyy0oeKyb4WTOH2oH4Fn9PgmDsdCAf3SCD9v6WkT
WSVCZBMXDJv1uyLZCFRml8x+1X9wN6tkmNuYOow3YjWcFAPJL8fXucuIrtNCrUrR9KzmOYfP3G9W
P1IZNtLhK28b4C9x9fcLz/1BxF7J3sidHBQ20Sx+gpSJ/HVcEL/8Dd7cfckSmA3z2B9rpltdqTDo
N6Q7a8FL6ljp2TzyLN6a/98ya9v36Nih99zA8HU/un3Db8IFVdVHTwM2mo/ozyLeLMI6LKQq2x61
iZPioJQbkCzo6CpLBGp4KWZ60ZPOpHy/5eeKT6a56RSRpxHndK8dmniNFrEDWKDB6WWuF7hXmmpn
/Lr8+5d+xgCSm8QEuBhRXJXcPoQTI/zqfdXNDLW2t9LwGZXOzz+oo3WWzr1hHDtQPZgBkZI41r+Y
8R3INf4zB7sTvAMR2qtR0ca4ZWeG1MZxcy3AMODNCor/bt+pgZr4RW8axRWfMk0Tufses3VSkb85
RJGjrcRZjS9fPxYlWD8RKlp1kkhO373krZSXwtXUDlJIt1lQ2I6y79e9H3xUdoMqbEDCrP09Zc9M
c76OUjiGwwB+LK9I+vLjjuUSpdY1Usl4qn9zTN5R7+1Kd/WgTJBaq7wBr9gBeWJ0cQs7SX96Eb6N
4CWMctdBjFQqCna9LILT4CaNWpImjmITEvxLVkXHS1NYc1oK3iTjNfHliojMOUo7XxynOoYG8/JG
cx0IF+6HqX7L9Ay/LeM2MF1Xv+eovv+jPMnUyKnkHziiuwgBqNCWEG//fdrhmKvM7jphdpdKm9Tu
Ks/Dq/WNezrh34juIgBs2pMNHnn4BgDoJoXHtXf0TVmR3pijg4WvI6CUQETeuyWBq/JkHzddvB0n
5s4W/Ib+A/JYQymJva8/oXrzftq3CZLx5ESsHub5JGrcS0qA6R5UYGLYIfhhO7btAzSltFBjgRQ9
cerYkuJyOXWhoaeLdWCeAaQX0ozxXsNzNPajEpzdRdwmVQNrfbquY+6E9plLzLD/kGTqvkmfDVsp
7EuQxiwQ5FTyOKm7LB83WJj2YPx0a0Nomz06xSx1N1Gz+h4HzrVM0j7gnwaaVD2c4Dlk66o4K4On
TNki1O/bf9uZg4BzVqyZkxhhOHTEYSJaGsoMApDnHrTB1TTSdnlo9okoQjTsiyukGxPGgib7xG2e
YzGzYefHeNrecn/0NJd5alhOMmLyKad6JtNamdDrMp8Kf9bDYSj2ndFIDqF86MoV6UWBxPC+EjWF
CVEBekTr2kxQH6wkaHxrWJJgV1mStgL+zSx/wYiE8JE49cLYcDYP3FxX4aKpn7UPfOzQ8j1ZWW0R
Z6JKLwn03rTgDAYCS3UYjDd41PBiggSjRhnlhjAvyjdMjlb3u2RXblqNgJWmVYJd2XPjUHsE+FZb
qJU5CWj5O0J3SuS4bWYbSbpAuZBVIWGGo1fZv8eU/gmSbdlpQmWGtJ8E7bLymBtowwLBsGT7mrrn
OzBCd3xy/Zp8mbHEGdQ3zsmPNnXAst6LWNN/5oHtQIFyymIHIbnQTEz84lzctnw31goK2TReTnUp
BgVRq71vBTp+S1ITSIl5yTfc6620JPq5yNm156DyCE4VcaksegPAQ+GqD++oG/ehF+xY0b9nCe+r
Ups04qLsytxs+7G2AfWpFG0YnRRLG9gIZkRmyB4FWJHumaSi42Hv6NrvfNyS1L0OjHbTed78kW8i
ogivsDA9rQPTA9wwSLEP2xGB2OkToWe5XVyXkSKekTSFWrkVIJx6j0X0brtydmpfYnqxKlW+Onfo
Dw/w9J/LSAEGTzhnESYefy3wGpKuzxshuMA/JaIWh7Z3DfP3187q16fg8gRD1WC48/YP4XtyfAcV
EUHwFoOQCoV+2k5TyoaGVhSKq/glrGSYicSZ3TJGUlNbTFknYB0CHp/WZlupuFcfeXeOKZ4SkzGf
5U+1gTFLxNK8/gygr5iN38beo4uhimSaT5asM//UcQUyyOwUIVnv0hJSNfTQVk0UTUniM17s9QUn
zd+idrmIFHF6+QeRv/AzxD6uzZUFr0NmdTOcX3WaVgkBKQSY/34Dvgq++dyDiPrwwP2VnbR8kn7G
03JmlHWFMb/VdZIFms6UIp4NkfD946cPyrHIxlrNOimt5K991U19/ucPRmXiao/A3VqQrXkxF6pL
lYJpXS6UO1cKPar3tX0MrCleWGHsYGhH2FvraI8qah3QIGXkJX0kp0EwiEv6zKntbekyyIk5Vv1+
UbFMc+y7GS60gDE1x9xkgxbZbL1ZRdi1auo1synafAM2jA84rqysJWqq7UqSkHlD87o5ifn2JxwN
xHnf4FipjVx/ZBghSwWIEz5FNn6sYoO9XA79yfpvY5svd8RxTwdF7IAkBbS+mzTvkGVga58sPiW/
LVjnTvHU2aRCIUJG4Adft4keQJoJevS152WwUHu9HZbs/ZUXvpTZPWWZ/0yoooXq7fXGJUIa/Kn6
N6hWGSk1SLq8a82iM98eEimGwAplHHV6t9HJgtHiO+7cuIsu67mgkqhYDalSx3n7tiYOdA0NRlch
xA0oK1lJMIxHLxYHuXgFsQf7nZCkA1LdV6D8OD/fjn+pAwUKrh0wtsQOiKDeko3Pl6nsLIllGWx4
A5V8cyESPgufpM3q66OTjhM9/ChWGoXkUIwY27v7kmHrOtQxEEbzVt67gZvNUyPgaYKa34zcMUUK
ITs0hTVRsK1x0v0aHCEv6XI5XO4PWCHPL8dtaGe0Q/yMYMgWMtA8TCDvySGtKQGCOTT7kzepcrL2
osB1rzHH7bzSp0qt8nIDEUuhWlQCBmFGIbrZJF+tMIP7WuSikb5N0ilI5slq5X6CfVVCe//houP1
vVET2EWR7weZJ30buhqguKbrg8d+5bzz4ynLPXBHJ75APzdo7NVhaaC1VJ01wkDBQkXgwCfCmB4n
AfPkrrxGyAZUL3631Yp5z1LH2JywvvvXrjjC/VUP6ePGSi4Ss+frOO6/2kxGZjZo+DQQB5l6nX8K
FptxqJoaQ6AprNEa54QoLnF2q/igHk4pcPYR5g836ZKhI1trow+TlcwCBwPr7Pc6Pep0n/n0fDia
y18n7DK6yVEe7AqH86I1PSfNX5pxZYNP6TrQc39/qS99ycvucW9Pol5PwqlF4FOQUzI8/xIWi+wN
PKudSsgIPAFouCUK/o6Swn2n/vSQLbGkUjnpxyf9iWESDfTECLj7dmqB55mFJETfIq47xkProlGV
7nrSpm53SZzas3Si6Gbz5EWaFTCQT1lE67P2YicEJWZ/L6pMSpbLR3VvUZ2u1Q/a7UIxSurK7E4a
J1WkVV+/Lf1gwKtAyhEIqKrJgu/8Uor1wCy4fkf1dzn0YQDU/ePndGwEVcVwQ0rqcdMqAZuckKpC
CsHM6/+EvMCefLMg5migSY2kibyUAU7OOkHgQCVFgt3kG6OpWgkEvEAj8gleOz/cklBD2xDUYMtV
4fM6/LR6Brn/LMNPFMPXxxuQes4upH0sSe7CFvnvTN0MacOZhb2DAt668TudyhOCVTRUKmDfU0K+
Z2XvCDOtOWbW1Lb6JiTdD/RASbSH4wtyBTUjCJ5LO7dnu26T4rExwfUd3gJrBzSKE2RUUNqAI1g8
EmWWw7v9NJGpVcR7Az/8AcoIeS+NSQtbKnwc6d81SMG1qXKkCrE17tzvEsp9gjG1OH51+C3hiJ0I
p3kgGZJHQD8AwjdZ65Anjd+ryfG3lHrXOc4moEg5IXKlLC6Ywg8qW7lPn1ZjmE8udBJ+hr/r++IE
vuNST3k3nw9iQrYhWGjRQmHUHaacxr1gCdMokDn0lFFXK3em/qS2GfZMCspim0YkRV7HbtdVyajO
KOmNYVAdAjrkgPMh7mbjIY0zBq5U/f9ftGmrbjHOurZSgaLPSYgzU9Cor0SAYssYNJZ7Enl4kwac
uFsyBTuS97kCeCPWvwFYqf7/bFbA1OtZhczpO+q76D+4mx9woZwGTJ7kAfj7vGG1FX8536s0enrN
QQkcVJjZiZsyZde4zZI0FO2rgaB1n/mk9f8WPiqZfJ3yLAJETFkBHYuv9h+/PsjfdFqQrsvnPkSW
Pa1tnx2Jd+g0ZLPVKqFYTPMOtMo6yKlYhU2S4SjjVxx41xUET3vnB2QZMLsdrqgVd2lsNNrAntpO
9pXYjejUt79Pv1sfuaPDzFWAVEqtfylvKajlxBB5Jn1TOv3mPyA69Ls8DIKbnIEhNl59RK8xqqTl
yxs6ATj6Rj+xJ7m4lUCcIxgoitVOiiiJDkDZ0dJ+e5QHTHKWAAUQor9csk6VBCaEj4mtc4T38UJJ
gsZwksTZYto5rIW3hTfTRsn3ooGMsm0ujG1OdDoHLv3kJKV/JssoW8b3bM+Xl97tMdKZW2lK5Lq3
K0EpaSnAtJ7nCnPrrdK4PreZ7Myue1k71VmwdKglAp6da9KNMgB5HXHGSTvjNNaTaruJi4R2a4HJ
jr8XVhGA8YprySWhqdkfu1Xspmy7BL44NhVjFf96goIiOJzHhZijgp82xFNAIbrNJbRzzGnIh4oJ
CI+YSbR/xuxLgSsS1KRNHTeSWY3dSe3p9bSUiC7anxOO/CDpMeKTeW2Qtqa/atDUFnPziS6yhNWt
4UT/NrNW9FzsNG8eCXDkI1Cbaeii/HDjpKUJLoMPhicORQgyMwDBUKXXdhcZxNGs1xF0ReJ7yxbd
mWOykmgL7kPdQ7DItlyTiLxT8Qum8T3qG5HZUNX3oCzoA7iSsKYBRijSfXxJpWjhf+22+90mc6vI
aELrb0k+oRFJTkEogtwB+AlGH6Qng4JHW4xF2pWRitz0Z6y7p1pWXLZoC9U5KqbPV7/XPa2cpaMU
qLU8CkUhU23HWuXCU67gHZuiJ6Ns06fWdWydzcsrLFh+PF25cF202OLbVFCaTanrOYUS4jplKyVx
bNLgHxE40UZPKrjGIh1Wv9LlZsSUIFEkDSztLEMFLiNvUOrijQKNUCk+FPIiCRbJ8zml+XaVPFMc
N43vvf51T0SN7vgT21amdMbkH8ngONemzreMVLHWqPOS2xA64Kfgd7CEuTGN1dKr5Jkx7MoLKSBL
vIkt6ACLGHO+wIC40YK19FqgCF94uBviMUHWqZCfOyZHo+pYax0ejFkTjoQGoSc3KHuOPEj6u8ZB
sO8GSYovHftPM5XNQezSfW2W4stUNpSFK37ezn6zmt3IBd0usVJ8J4PA9lJwz0Be55KfKfnmlHzh
7V6W9ELyovaFymbfZVLHOCjGMJ2imXlXtqwMVPn7XnmgMzR+6X3qI2cVNeTxky164XE4peUoMC4u
AhiJeLmuWu64JzD+Ttt+VdEX7+T0GOqEc1KqPkS+JgbTrRoRfIHaTNr4MqlOtw6d3YyT6EaCwFda
BJcH9N+QVYhU8QCB1xfqC+jhSi1Dto0OKFBMMxHmwHHpxEGRKIqWjK1j1juc9yBr9/jZsq6Bjbs/
RIfQTaF+Z812KaIXHHu6MDZz41FEydiZYiOP1Jxm+sGfdY7awCFV6rwr/4MQ993msRRW0raXlq8l
zbAHRPsHcUvNjkGXxnoAP05kAGf2F457EZsuHkmLvbGVpZn2qfoMZYhTrjwtO6DGFn9PlYbKo4i0
Jvr936YZvnxMjrU80o3Qnu62Qz0Z7YNnqah4+5t2ntosGj2it0uQvAUcukurA8tiqV9ewM8RElMG
fNOD2WkuRqxbKAnPfPmEyFbakkDbqKX5v8/gbBhz5loALyfzMqQ+VdlZo/PauuYjuoz7PKhsgYym
YyOMztdxzKr7MYUjzfg0iqWyg6LeaObn8UDi4eIh84YtfuJv0111ryHaPnFQgyCUY5MagGTIM3Z8
KPQWLN+Eqo7WpAHrXyc5oiPyAdlLd9KdRmsZ2H6v7qk3V+A3jdfUwWmJZfsCAWCPblWqEhx9fgcj
zmXprvzPs3emxRShigym9DcWYIle9fnoZnx32L+TXSv1cnkLyR69KmLEvZ3f791rAxQYolY4/GDR
oWf3gZXFDhFagZT26TzlIWoT96uCTXWFGAMxjGOzGUlOO10MqYJiRjkrxwvyQbNkM7rHLqKyzXSW
sV4yFd15Jm38ndnipd/l49wcfpviWEFl2Y+YoGkhg6hPcmhl7MZFnRO9ItcDgWSKo/LRHlrWxBkB
2hIvr0uQh+GC1V0o/5e3p//Wrug3oBy6+i8ZCx4j/WDHH/fM3w8puW5i//NPp0ZeL8w6AosQpjks
xdEq8sgmemo5qpzrHw3kv0s0csncaebiG5HKB2xwyVABivGkUQhBpTkWkIpFO8y98ddWFcS6SXpK
KBV0t9vU2g+q6+kB4uMPuS1nfJ1Vzrn8yyR2ykscg09CfJ91H1z72SEN+NxCvPnZCO95e0qmqBGe
FsAp0Bjt86uZgkWPItSHPhU6sqBiCzPo+V83WVxAI6mlbK491ufDk96bZwTonZG+KkaKBtGE1xD0
9YrDu7/OCt9NPvd1OKFVbCi184ewYICBETz3/z2eDyOB7hSDtpJOFp9t2GJTFOhShYsh/HBs5QUy
E0Xo0qYVcfyiuO5dMxxMS94D3njiUqU5TLw2keyCla+rXlBMOCKIIdnVJU0dgnnw4cgHnprMfOc7
W60T8wV5ZUUcmNj4gmCRn7k3Gn8yYbQRYozoAQ4rsXmkn8Y3miJJvcG/WDuzFEQJ4hqhV4SN1ABi
4+G0cCxpsxNWyPis+FYKvAXOSUjzSwjjAPE6gjMvo0+OXnjW6Gknr9juS9QwsbVC/S7aFG410Q8E
GuvDfbbucOMopOO70++3l/W23nxaWT+E8PEh3g63epuGJRs9Z4cdxo+pOYJCBs0OPK/McGZuiFt7
bpySEKAnJcjLycWfw5YtCFz+se5YxxL/P3PL0/yld2DF/Ey9YzSL79tiAk8wTbfOG1Dmde1s222F
FV4oNRIVZb/vUNZoBRwvY45qUdLymy7+2er0gAEqH5tHDzOQNUg4PKUCFCgjofNpEkZ9PlGjEez/
noknxinhxjXvpJhZshzKfylc2Y3nn83/8phacGh3rm8XOu63M2GYvDZi5v3ce+nIVlPBvCKH4spQ
AHvERDVkpbK2AD18QYRwjtk4bd1msB29mIr2ZG+FRQad5/Cx5W7yzmgDIbENxpFrgy37RztHHARA
RV8TKZlfDbV/8psDjeKWhjQ74h02bxDxPpnN+YDDVbLfHfKjeYTU/BhDQtLhAg+ef8cJtjKZAePk
S8Z/bo7xHnIr9e44iH7ngt9gB9pycCh/FW+5kYMY5Hb0QsTPnTTjkUcULEqhtWuWf8u8Jr7tVkvH
Nf3U/shaVrFBLIuCuQWCOk83GbMT2Xb1+QlgfrPBgLSIFrOgCao/KG0Z/lcnt9KwvqL65NeCxWVS
80VhcZbVDTsrlD95N1R9c8/RkqQeRbnGx8DIh4uvuy6WLBL3c+l/Y2yLYMjf+hyu3u+gLbigj5tP
LPoHaDca5hnEYxuruH0pHSKLiXZpw0uxN9KTXK5nqdgP1Yfg0DyAwbNrXycPZ4FLik7Ly7VqjkSJ
J1Wunz9bSa0846GqCNZytuapoaYdgt7Cq9MpOUJ1E0AiXioGnNCQtzomjJlchv+XfihWAf2BSBE1
NWAvas/9VW60eavR7sE3Rks8uwVnpr8aVFGSp49+pviO29xNvTJiUUh0fqm7BeaMO/utXBFkqPKe
w92aTIiFTO7O1/SyTtTl7SDN+WLd8FKSWGoCr1DqRStnVfvVJkzZ0gDG2nL8aDkr58gM7uzKmxLY
qmpRTTPlmmwvP4vydWxq1wtfiFt2IWRncsFnTpkXNsTcAfCFySHh0GCRpyPT/kIUqylUVqfjzYn2
fhWU+P64qU3bs4s2mZoe/KYtl/PhT6zXme6odfrytlx7PG5gRUdAgdT6+GHNTPl2hT3v/SPp6xDj
rHmEMDUaukM1MdgbALO/6QD+7Ufc96fXTp5OzQt/alvagezihMae1WI4Ilz7ENmSYI7YBbLY6o5w
vfleQFku2adg63SXYbdVssNEKH3IZ8e+sri3qQDNjo5LvDea4pdAULvQgSLijJhp4aC4hnNjO8oW
pmFuH9sRy/uhiGFbYWQjBrXrh0tqv620BH+Gc5jpv0yquIXG/pHJ48jFbNEM5NGLiNRkoWR7Qz7H
9riHW1tKUHh00i3I3EhlPcGm7bZ0j6TNuLrqdfTV16A5/hErjVQPZLaATJodGFjj79RRdgumb+Y8
uSJerl0eYnrBGoBUlAcnsISODGt385Uemvv0YeS4bT/NkCjlvv+ZKoxz84MkZchs5t19sPyMmHQl
I9/O3nUuCwcc9z+jy4EDx8/fWa8CSq2Ggrd1tLng9l0KlM8chaqavoI6qAyTAMj4O70sv24QoiJN
MDHqpFV9rFKKSVLL7NkjtPX8WCzhVmqsN4ZBRaxqBIiS1g0u249po7AdHyC/peuEgZdf8SQFQpN4
RrkfIseYq7df1i+QhF6wyZ2Gk8QCPAZqMGn7z0/Pg1R1rywa9xAI5UzwmhIdDCWnF7qcGAA4DpC3
elcPN2Ej7tFj6VfqUSB3oRjQ98p+ORf4oXkNeVkLldm/QjUB8f4NmUSiH6LKYhEYHwQg7Ve7rO0D
kckUj8Jh/djeNF+t1s1e/Idfqx3k9GuLnRQ6an79hSbxm7IvBDoQvXZWVbUdPhJpRZR96rzEqi5E
AFCC3qMmNB2h4tQsJAS0WOpkf0MPp3LXEKyCZl4NVluFq3YJg7rjj2GKQ8FHMdwWYxf4sPz55Ace
StJedUuSaCmzI0RL0B3jhiFxkp2KdUAxmriTwIXXFuwWE0mKkYV86PA46N2Y8ZCZrtvyV3hOOfV2
rdTRwGtSShJ84XPqI4d8pmRlfsZuZ7eZvDciwjzbpCTKarCp00hqWyV70YRxnk4JVdZQf15V/wRb
MCDJnMS5KGnuZtcHNOVRUqSiavELHHhpsK8hQVRoyIBMdYD8wwflaJ2GSXJDVCiiIuS1SC38NkaC
xJNUOzwt7mdgLJ3j2dv4S4867MB15ya3dkl/SP5+RgjPHQV7Vg8ve3u7nXGmw3tj+p7jjKnHrN51
IC5+rR3fK/fZ/9MAx4LgEeiEg0HHOah5JCxYb1AF1vrknc5U076+MZeXMh0cVKq3q6UpNVlUO4vF
KSjW/a9gp9kdhTDQDkc/sa7/0yiv2SwYimw78sz0esoWPR9O6Ri81ZCvDgXK+HKX925m1FKq1PAf
urcOVhsJ7HSxBSHTY+8Zulj5luumKnrfBWiA05tfA06hCCJlU+1I2Flja6YU9V5ItqyEl73kFgXQ
WqbTDaOuiLujy2Sw3cL90wh8N4y8H7KGYnfnVFR3bDdqz7A1jrlhQq2txsRsiCLll2cIulp6CmoO
jpIsZy2v2SreH7n9wq5W6GU6g+KnjwYHatta19wOZEoxR8+es7XgRZEZNc1ncMvGHMTc1b4p1Bg4
tl/ON/z8N4781HhofZEMl2E+wXtuFSQj28rpDUgIyQ5uXH2Ys4QCTI/c2nKxl+Rp8X0FjdSXlcYA
Lap7f2KsS5M3wWqWdUwL0JD6/IRn4THFAIQ3teoaxRP6oY43QpzTwuyTUTU7JxrYj/iWlkGfSgcc
n5e3iTtppSH9vsSEwSV3H0sPrc/RNUJCtYx0sTHuJ1vgVlLloF2bqIrT4hR9Bz6bafSO5ahBxiQM
MMTYGcS4QXAWZX7S8LlfnpcKkt8EGiLPOX6bzaIgKOcIuswlE+CF5hVw/dDE9bgaw6CltfD1W3h+
w1eZy3+UaB/rum3FAuXRe511qNhZ5MWKbnaS+4/YB/O8uOlo3o+DVSIMjOwKJpzvQLaKpi3WvAG7
9NSRj2Mmg9+u8SXIyPc43mfPSe68sNL+HHnHSCR19MofulGXOrk+3TCYg8OFbS70A0tAINX562PN
uy+EjpCGcSD2s/nhJLEH/qcnsJq5bkif03N5Um9Ogw3wVxRNPupDMOKilHTqox8gVNUK/xzKhpDM
Xf6f91zogcgrOT/RWJhFTp96X/69w4QnlDnfg4GjsoIVg1ueMCiMtER6Rpl+9ISkVbkJcxtSC5aU
6sW4wrW5gm2hZIyMxgyHxhDQHLUVr6dD2dcSekLN64S78SZqC8CcLJ7Pd3+alom45hjbhqm5UcT+
Zheh2GN3iSg0urRaTcGJgKfMBWJAdhyj9J0imbCzX1Ooc9ZeT2WprrHZW9VV8xFtqqhXvIjdfV7v
rvVYyNhZXhkfr3Hq8rQAIVV3JFXoK7K/DG7o/+tFaigcfuY/WIZbvMc1RbG4Sfvduyq8tzUV9ckR
zSDC7eK1VFVf4t5U42tWGzwND8lKXJZQWvN8lxhkQfZjLkcxGfFkek6FdAUaENDIIFVpeqofVG/6
bOSV0T4yjMlFpMUhK+ZQyQO6T9D5NIQfTMobLtMccnZKF2i1R7D4I1gxyqdkxO7W5ZLuvIUIbAjW
lb+D1kOUcITKmQ61/MPfr50xWQ/w7Dm8IDafnYZEVo3blVDqKZCL2LuIWB873JzaRIMlQMA3hboW
GNfgIGhzPRfqcJ3n9tk/OB/wCkwImLO8rG4EzPdVTa+AC5D0g9NE0eLidv5aBdaNXxM/3rRl675j
sTep47FTW+lhs+u7Fb91T+7w6Pnt9P8U90SG3ohUdRuzGA+UR48OkiMAsncVxKtPKrDgsMNJg9NU
TinE32AUk89fGe3Pr+AYouwbsTtFru3FS7TDZI8QURVyuwYxEeJnkD/ptbWt1cpb2FjehwQaREL7
MgJxLm13T4VqomBOP4iX+KqzmmWQ0b/Tov5yJYdskGQuwEOANqu7+tx5rMV2fD6uJbiQjfPu+REm
Q9baEZhlkk6DQdscXQ6AVpISDsZnO79kZBrtAx+xc9B0eQkAQSkHF8XM3YyNQMn1J0mcws2pRVny
rp4N6dgNl1aIU+LNC7Q7XzO5HMhTe539UegD/D3TIRA/7gHpuPaqiTbjDcJM5iaHSmJULwZgZyFw
oyGeePGvLkPBpaC4eDAw81UTD9uMUrrgafHlXV1u/3utpnSF10KqIkyoEWvU8gHr/WL+akn2REr4
FUF3jjXXc8VQl4jlw78MJWmzMGobuMZ1HZxvEHmFltQkybk2Qo0i83hHRt/f6y++l1FiWEFQmRrq
69VSUVL7HQEYqKVw3YF/63twCwNdpVJGLOl/18XKn0+KGxDA15y7UhDx6UMdBgOIZptfc+hegakS
A01TEs3jkiKazP/s8D/1XnKrYXSzpZ89ypgypjXd37ckMsAJ4o6TqKu7ZPtq/2oEd1YzVvC7TLTk
D32QaTdwVVP7T5h/kbkqjc5jsQU/6TVgEUBPPlfNokHjaqFX3lroJQer6+o8Dtp956fEt/BQOHAc
DjdI0O9DCslhKXkMkf4lB/pJa30thqYrk0tDVHfKx2II4ZUIrwm++eTt2GduqCTx0f83PV6ZnrgY
6bHMa5xK/iTVfLjgRldnlp5a4qkVIhr5S3Ue4Gmbxpvol8negoe9N3Iq4GrCEvTkDuH7WHDThauA
58FmmtibXaG7qxbeBemb42vmRW4db4jt3EhKaUWYPQ1G3Qg43Ua7VqpKZkGMOZzZuTi4hmJHHX7h
5I1P0UPgqiauupfjVBXlLQMQ/HgXCQaHQ6VSTisbc33ZxF6c7CWukxEBgSWg628BnkiStLwqtHlP
gX1m6EsWb/wrok6SL1TbukBEO0dQaUi/EUHKZ5nNszI1hzfzLPKZU9eofDM5ofBBzWB1xpSDLJkL
QFvLNZCHgQEjF+t0AYg67MeLLtoJgYN/fyoL72Rj3+4tEu5XJQCFH5az8BQzWq9/tmQciVd7qgJF
NyBTY+SYMxMFoS3yurWnREAwmg4e733XU0KZM/rPmYD/BtybZSrK0PxrUeua7zDIeBZjU+V5osGM
A66nwJf1TLSzJvIZs27HaTs1fD1D0k4rK7gBY4+p8atymG9y30cnu4VGAPoqxS0Q+rICZeyMDOYR
Zyj+otMTrm7s+X1dOIz0VPPCkdSC8AXQrA+EqIInRVb7qPVPwTkQk3ey89J3YBo3BckTWCuGYFrJ
xB3yKteRN0obdFrIzSfr6cXI9Dpu7+iAkBHvqBe/q5+oPqwPYdY3xm/CE3cw0PWuDUDtUrgw7PsY
+f3DQjfMftEDQ9uvzW4s0JK9UXJF1faw4sFtX4gb4MuXA7oCxpXtOCK5DoDVC2RaJxwgBgFklqXB
0co10ajMiBqHOu5Rrhb95jHMEnAGh3Ca+ZzyiI/ZW5/2xTVBYvmJ2HswS8H+ix6ob5Z+OnpKjLFI
zuo8K/jSvjlrJ4PD7ibv2l/HFw86jPGfZsJcpidLaMaYaWQrL+5tyIH5UfrDQVZ4BfwRWRY1iTqZ
oM+pBBUkOajKayLTRRlqtsSq2DlMinMZnlhh/RtCfHUmBkfCeC97htvZoIL0jl7qhJhv2Yl+PZUt
GY2mK/ixrrdRfS9+BgL/fp90Ikb8Er9g5maqor6nDU8uAmA3Y8QGc6K86WhUf/80jbF/MtgCcjM3
Lpc4l2VVc76CX9xeaTqFm45V/W/L0q4QNFknMWAx7MtwmC69UFTMCnA87yribW3YDUhnItrF+zol
Ba1R3oafayONDW3wTo7Hz39xn6+6A/cvBQZtLB3D6/dKi9YyAyCwJ20hrX2JIuI9eVNe8G8LMHDk
qE+LkVO0S4jc23IKg/En+VPr3/6kIX7AIq2nFL+y06Q63LN8oOkRNCH5UJMVCsYmY13QwSy7M+Gf
aALCkpRsk7wdrB4kzZVEgxgL0dB6LsO6fRxN3jFLdGYBtNqiZhq9gyM7ssViGTX2+qSQWVxxCqr9
voAKYgIKZoHELjnIt0CvQ8XIakxhNHMp4H/4BzccCC81XYtFt66RXHkkPdGEoPUV00f59OyYPO8T
6RoF2rEVeh/JeH8HF2bvjKpsYhFI/99tB7I9qLY7t8zEGoWLvnrDnJNUR+usgHJioBTUV/DUOha4
1YRSVTO2ZL7Jl3lfALNcfQN+E1Tts6USLPjjFfcIRnJS5wsAYvkLL6EZh5Vuuvv3n1T/7MrHMJxq
7CCKjQVDI2sTtbR+FxNTyAmAMP3O+xhrfJhiZIHq0ECcBLFCdes55FflOmHCcB/uH4eNLJpyZTOP
KnYLbHu/uk6HeHaSOO7D+WnT1yXiCpMKR9iMfs/P6J/aG72IWr47A7na/FWr0XX7vfjj4EADyVVT
jMEObH2Qs9/gHDDLngSbgGAW6tzCfJPIf6M7Hr7ZCjaKLwugNYDDYaxIi0WVN1RYrTFvRk+636WR
3CYSxydpi+BAJ8ULDf/Qtv9fU3aEE2lIbkqTl8bgB3QouVxvgui2elbKerFpAYWkWat20Fma9AfW
PQlMSERHbeyApKgxk81jlx2JDo35+5BH2bqXjS+YE9lqUHdrm5AS0NiZhZrgJ/qHHh3UZP41Nqsl
xrtBmJO00HtNvbtR+46jwzo8DFgLmkWyXXZXAVlTwS78ZR+mifaFMUm/xOBQgenlk1DRxO6hJ6Iu
T5IB5ZoNjFNIcJspjRabVerViQY/0WhhJxBaDe6O1yLb8XfUnHGi87uRy5qhRCvAvtV/bEo9aVjd
dJnCautnqofmqt9LTy1LJmtiETpnDJ2vW06cmgJRWm0C3ey+YXHQlIOnP8nwqCNTXESlo7J8DCC4
W2Yfm1X+cjtRTb6XfI+E4Gz18Nkng//RytGfd/l+amvYXlUseJn7mdTNoZD+uwM3qbUbOTLrMFzW
E72/qvMIbgBa1SSDV8MlS/kD+7r15nrfb9DER/SXMacka8nX0jy0qeWrYEIr98z6CkDAVzRJ1+8u
qTWsUp/1tKm3ihSgBWbg9HzYxo7u6mMCTezA7jL8cCXE/xOGeTGGRLi3hvZZLq6ybZSOZ6w8AwKp
xQaEWvzpe3Z2ZIuNZxTLFqfQ3ny9+oEhEjCdar88/M94Xodxwv9jhjz1ZnGuHM9ycqFN5s2Co/Qt
dnacilrA8PhGe3lLxWbL3kw7hrmnEoxz35OV/rJA0JngwfN9wxrVik6p5SUuwqxrn8fsvTnhs9Fx
5Kk5C7EYkOL2cEXvUFISq7qKUv2wytqIjUaxLs6b4KzPKv0h7+L9LCVzM8og0fIjV7QlK8b7t+oL
WC5wAd4UsrQU/wJUgS4DdxCrQOv55mP/Sj7s/YPIndhnjGsUNlmzUkeCQCtl6ooz2gbNPXQkqhFp
mT3zHHu96NmyL40l+PY3k6YkhnvHafmzZHxAxhXykpe0dXTp2hGiCB2POlGL7xwxAY0K9AR7/s4i
AJwK3wg8C12Ff9HVfymNpY1OdKy/UAb4cnZ1S+tlbA1F80zkxFZrioXQG+PJUMDc9niYUdAYsNwU
BmrlykJSSxvXD6T/louLPyt/cZgbIgaoWUFLYsWGfSD2dVZ0pT9QZFjqRDSa5lEAYFu7XYK8LTu0
v/UfGv8sOE6Mt0SlJGmCrhVDz+/i0JywmincPEfkvCuRwmjGDDIet4d/w6J3XIHD4KajUeZ0N9Kk
OSnFo7G2S8MgNyxJ+QcN/8i+Y2OdXbllSFZ7CYhyCMgxEqf47E24tY9wFaige3CbI33CEqpi4aJI
QDFnXTp77qtt2KhemLsTlBe/ZGog0GRLN4xUbak39XfNCoUmoh2+ZVw55JV3FYC9O/uLY0Oo1PQQ
DGd2DnBbWXJajYpG2lIa+7g26P5b/13p7k5jevVrP1QVKDuJ7QruSvV/g4T7NXGzBHfMsY12N/FQ
utwZSrSbb05bc8VzAWjFxQAYjHLQkjWHmQ6lOhZiNNVeQ8FlLRy8SEhnWHASvDcaEmFiOWCK0O4q
0frKzqObiB3yrveJmKfc0AcViZHRSDdILPYBLPBZOaXC/SMWfqkr+Rs61QbBGOQoUIysTXBY9TIa
NbTPMgIWLbGA1Z44KneYdfU5W9FM61VOX9ZGGbKUAdxmHBM7oZcGGli1ZYLsRVZqlOGP3U34hIIT
Z7ie7ZSE+JJuGdsuUqcZ1iyTl+svgwcc0raVsyYOH+UsVZXZvdbpoVkmMg1+y2eM2melEmXA8LFa
yad1dbIFQ7sY+v+3j3to0jYupJ8PZ0IS/ZLoKUvRve3ulyVsvCJIPPsKFNUfouVuEq4enGFczJQA
1GQXsv8aT7wCr2XQ5uVr5dJM1t6G+3uSqrBuYJ39WUE6Icy4N9E0iMxwzK/hF6T0X+jxvbp+ni5W
9UuGO/cBCg7xRenzb0WgyLaS4JPAxvPOjdHgDC+X6e96CKGZRfrn9djWkWt1S9IWRAkj049gBmSo
u6N9OoBgc/LPKNJazIVGDW9qnXdXC5NdGUwhp6MmscFh2dt2JOGLzCVoAHCY+o9CJ5YnqWUyh3Py
dkUrscSDhv++XsUC3yJQrliyG66QFNDjbOzec0uBcc2k86TFqoPCq5CVft2byuPsklSSdMrUmz/R
tAjsHrCLm5uPH+fRs/eA7B9mDXGkatiuZFATGtCru/rmPLaZpsiMwqFgygFmPsYPjmGDnxXYswoH
uDUWlL3ZF2wJGgqp/Go0KoLk6bz/8LsVZaD7H6D5Q9mB9BIQTKxod9wrm9VadNA1hVO/rEg02t4K
AtY4kRW07kP9zQK7YVdaq/QeIgH0m6bh4MC/89ixGoRE5UUtJ7GMwssecKO4XqtmV87a/j34zNPl
KC8MaxpnFvr6a1JIiiVMeg25PaWUsdLQqFd1wWfT82iUV3LBkpdqcwmpGSCZpAxLMPBfzLJPUbMV
9NY/++3g4Z0cqDCFisAcFsb0e7SJQzPF60iaPTciciadtUEukme0mXqbhndxUdM/otztLCLnCKki
KVioLB/fR2okH9RXsgckXMJp87GDbnYLzB2ZF+lWWT85mBgFIgGlIbgXntHChi4gjM4hxW3H5S36
dWT1Yr7O8LrhYiSDWosiBq8AHrUgAQH8KNaZTEg2eeP+GVdxYWpqDpUsUsBprKDzLbOf5CRX60Ty
dGha8nsDTIRrXJj8XTTzfmO5vvyRTTWO9ptc270jRMyXuPSdL2qfVMKJ00Ce5EklZqKBOx/Iol4D
0bvYuF7f/ZMgQB46KJEGDGGOStE3J8aFbcPCnmRHbswOk0gCyHF6+bp4Z+5gAHrqMbqz/LItjvLy
nd7HegJ+mo2oBfiopBIGt6t8U1sgaqrAcxyIHzoX1vOQj2BQmwZYeFTBcFeR2Ts0cgq3Efrx7LxW
8KkitPOh8jTs79aAj7lAlSGbyLLaWqqSQ7Lf/sGfzkFxQZ4eV3qreSUoebhBSeUCaQkBn269rTiI
k6EG+JI6bEeUtgo6kiuhilAJqblAqUdnI6SKAEzcpMmZCBji43o+u/1h4/tZW9V8I3uZCzyCUTSI
9bTpw2tTFkBeMPrEsJHb0EXcCVK0l+MFCJBTBSPO3CqYYXDWmOEHdEC0/VGPyw8hFmf6AGoqmjtN
6anoU77/jZq2cqgOIDkRwhVXjNMWRAS4zkSlwzEldvK7l1Qq1f1ZA1gaTmT+4IYTh6TXPPzST0HN
kxI8ag6O6rbG418Gae9O+DGeanfls4DyK3odKerkKRBQTRgl/KJPzMXU8Qrzjm5DfE4dNNaLIOOz
jPaKoDs/FHcM+Sa0AITKabUthPra7r2CJz0y7+gqYXd87Q10Sk+3Mb+s8nZMUY6XQX/zwfcc7PuP
i6s9SA8rP+IOYmqwt9Of1AyReSAM95tRnaAwWoZtV31ME4cmIIDWaqGGe07QBVVJOy+2POPZY6Jz
drVLyjetmqGuopM6MAShF6ucO2eR0O21fCHJ0cxAfsdiRUg5vITi41xR4J00EhH73pWV/jeHkKOL
IEFOF86dpcLzszzVrby16MS3HDLyf7svnbn8NtCwE627Wyic6GQTMmfgLwqDoBwg3pbXitM+1CG9
gc9dgagHr2P+ogU9rqDjLhOHSuep2bmzpbP/MtCndga0Z5S4/Mf4XUk33ykUDOfKuz7hh0jO0D1t
H6BevHlKUhILTVQ3WXQ36VXQrbnhg+kGIiE21+PvdqLKPajhs9mJ/18y559m8DW1DofNt9G6Rq9X
fhskiFApSbbI4S9+G6vESNIXwXRe+nkOvF08YQw0JVnk0HeFCuU1B+qxqd5qa318ISPiiyWyJAnq
QcLbos9fMe7EfBhnKKr+13Vu0M8Em5j+i7xcoN5D3RdH1HpIYNSmgXVUNYy9EvfpMbY4822zJyxD
mmfXmoFlk1+Ow+eGz2kj/vC7397UrymTDpV85WQU3qFnZcGtyacku4O2Y36VRKC4jqMJ27y7GI8b
oxzS99MiTCgQhw9oSWeD9KQDM7EatOHAe0CVJuYrxb/hM9jmFzP6jAxpuBeQ3BLsq9+9mNfa7weU
hOp+3CB8hvFPnIb8E0ki1KW/7v4Stytg28YgbimMW4LdMdT2QiICySefIZaWwRAO70Vz/WboeKE0
74JCXWKopKWtj3m8p9HjF3q9O22QSpj37hiHTQDajyH96UjyoAytCZ6M1j9JrjPkrTjDmfikmebK
U9GxXcO5Rjw4mUNyMk6hPJ66S4Le2cnQdHXPPGh8sgQkthRP3aPcLxuRejRrR54sC1RIVGslDs6E
P8gxnnmn/x6b3AGcAprKj4fnalKJ2eYQA4OI2oPSCxmiiyOtDnO43Dw8AARNdSInXtNcnQ+p6/NV
eXjqX0CimIQUp79qTdUqdkDXSwezsF+v6UdZbAIUGoc1YRwHJAb7jePCzCQsl6rJLzFNLRPimisu
pNmS4QIs/e1UwfoAbF0ZO4+89o8szpTXTIX+37iCJKhZLEpHtGa3CHPIVcGJz451Qow6H6Lyi0A3
c3uhA05DUL3NeqSeEntgfpQIf0Zyi2FM4uXEmvIjjG2baE2nweklY/I8F11frnHRj9tUBCN8Dzc8
FhKZLsdKm7HBZTWVP+IEt0QeJXx+2XlgVyLn+QR8w9J0A8sLpmZVI1HFoK/9RAtGxu4Bx2a+uq/x
8qOF0PYlzyamEwa5b5COyStyTPYPR3yVk4BHhZeMijye2AlV6wRqDLiYUZL6UGzi32hduufv/VYl
IsQEpzhW6kV7u+QhIAYncnZf0+frV4FY4vr3TTWxsNnaD2ZOXZwlaM2MX+m+Q/wkU5Z+enkDGdRX
GPkX1/B3Zu5N6UrWzrdrYVadnqGVk46tzoX2QI9oawslbkqRP7nOdd6zTZ/j7XkyiIUOjjeqSQT6
KnDYy7L+hGLzK9ybqoTDRULVhpwSVSFf5sesjrvGF4ZZXLGDGbXnECl4bCrJZbMv0BseY9faeZRv
8ANc35U3dahMPS8ucWQZQGwGNsXleHQUwSuxNJopeaYqLfBe4ZAGX5PCjsquemuJoMaQsaQDGEQ7
crv1IanMGOEMeRceqm42XPTZutlafxRN+4fWG7E80183/zZhvEH/o3w/XCp2bImL7UuJkQHhPzqm
gM5VLWAz2UeYHH3q3zamS0GB0b8ZhT/T3UjxKH31PKJGOugycK1RIhAAe1lHzHcePuTooF9KeSIW
UrR0y0xJUTK3U8WmAus81EnYPnrC7kp4bC86+h32BxI6fsLgzbxNGkcEtM2+brshu+xZaKhmhiNc
KPL2WB8QiLHX/tkhUoecSh0zj1xOBlYFnuXy0GZer4Y/+9oJn20OTzuKrB0p8L3K8AZoOl3F+Wig
TRkYX1aeTkUv+IC/sFi/ZZFRmRZ6A8d8cPJSDJFzltqah0KHvyjh22iv6E2VHTAL33zFFMmtqNOD
MEeE4wv0NekFBF8lVHTacIgyYyv5olx3fnXp/RsF6qdhZOYuy2WgR6TXW7X/4asusj0F/HgGJ3YK
H4jAuPAWuEt9XVkRP0yn97CpN5SgnXR4tSYDqFdzRdruNsNH+cKEMCJVPJMA+nqzds1VBxt6cFIM
dpIknUWCpSERa1SwZghp3flbis1INBr4MBsWb48fnX+5Yu+5VFk90OX/mrL779GwA48GLrhg7kUl
2UcQAU7C5PX5QeoSPogcjv2zUCqRouJ+Nwv7ow0Dk3gJF1JRnvbMXEcurYSfn9lHBzvkKnO2pJ5n
5Z2uPg8McOhfYUAEiC0O5bl0wp157/RApYiwJ99VDDV/cuC8dO74zxBhqYdpG4Fdx2+PDcH7eDud
zv6dEhSpAuKQCRHd/WPi7OxmrlODwuBmCZEuls06UOdPGErgMrGt/Q0hyHZ8bcUuQ0+Ndyje9eZg
WCgfYRTntofkot0SQXNLT9K2WNnVoioC8OhRo+pAsZgZv88sn/vQ20mfpSYqO/I+Jzd2ipdTEx2e
3/5wcDrqlRmsg3sF6WxnGeyIaYka7sLH2w5lAuSXmMhyDa/L/9dW99Qu0AOsujtMbzXB9mj6+d+f
uCqEk4YUS4cyLXXb1nqXRJaf3xQPa6fkcojJ8LztVwM5A87Cg2v93cKiKRHf3Zw7J24lWtyWUDU4
iYM6o41i7jX6P8VT+NLw9Lv573iOZIv5rnhLmqvimo9e0UlFf9Z7eOW+Ej8qAsJIk7cYnAWF6u3p
xByRd+Py14VC63DNYx+1Vb7sl+qtnECBztJ9bucYBDgB8pP8VrNKpGwmPJRk/iMhTNeCP4Ewd9Up
Z2KbkV8I6IYCYSJjlBSJqLcDDtqAH32HMXsrGotCVNGOtsumkQRDuvv43R6nqpvioyf5odwOVnnE
zbyEEoZTy6I3imE2KWXfP+HHMIl8hSfljg7lHNe2usFEDUFHvKEPitf2dKfmCo+rXT8ODPNI1QzC
SqzRZNnNGz4vwGWf53+RpRpvadgM5mPfduYIoItDJVq2sEPvSM5WHyNWrSnM3GcFHg4kAjjH9+o0
O7sO97K3pE3ADHm2KRRREEB4Ykyud+ra/V9vYfqN3mjF61o5duBXbs8ZZqZYz/uWGdJymy/HfrQy
DaYYoz/A275/tmEupoj+XTzjW4vqbQ+FzgMTF+U9Pc/kp2n9X0Ev8pD+DR7WyIF2udnXCqyGqjQI
C16liDepV8+ElUsXa6bvI6kgNflM3dNPeNxEAI4KtnwJh6hWu1Zg85xgIi0bDV+go23cbNWDPtMd
NTnZEr44iNG6fetGJQxNrUIJOIfhDP5YrTq4JkPnpajS3JMQAOkYO40+Q5O+XMAzwxRS6TuhnviD
S/2VVsOW8S0mpScujFw1oGMNg8b0Op6rOXMG96fO9tJ+N7zVFgOT00arprppy5N2H3PwjMtKCI0t
sM6fCXPOPxZb0RimYu17fWWwRfWuyLKu+yw5khzfjnacHyc+f/Dp8nfhiJh/helhph5qL2svogDV
raPoWJltx0jZDK/+WtOa/LbzqAQD/xAOiFNqQvu9y2Lo5pDjFp65RQdyxn6gpjLmy1LBriCpzNkM
xeSnmx8F9HJKmswVnU+8qYj0hitYsB4XhBMF/s5xaA6GREerJE/eBClXfKeXagxdKGuI/znVjoFX
MPvnjNYfNrwVy9NoMTRwE9z1bKe87tiS/bkZCvmYK7tZ2+Gqt6SciUAnwSzj7vu0Sn+EOv2WlvD0
rQVeP6G3ZQy9RWFgOo6lsWokOqb5DGDOiEUmnAu/tJuv/Qykh4vI0QyfBwUHmMrhyHULrQf36t26
D7XuBX4D3hLvDy7xJu0W2+bYo31LuPh0hOx06Ulhq5jaNU6ktSzHvqeuohbOb4NevHvrPnGSHdDk
zlvug+Ckby+EPN1abFMK/Xuk36k1VpsBrBNS9We3UrjiwjuyDxZcfAs23tZCx8CIaIymIFu6COsI
I0bhTfN0HuQKpr7eJlUkSuv7PO2DOtNYE+IB8B8/cP2tXsOsX3Q+WRhUHtw1TuQn+vUAeRkj62Z3
lAPkLlS31J0T+Y5Jdf2jIxhJrttiTL1UAvM1I6thhdhuH7MJQ3Y3O5sdegt4101HGdNW+etwLBmP
rjSe+DWBfly9nuFThkpvOx5jzJN1bG7J5eR/YZxAQXRm2pIsNxjMqnHcSEb+tHWtmliIlUKddv3m
ZMp5rIqlCN8G9AmtD0od5qjFJDmSqWkfqjCeColMiYUtiHyAsdWVkVhXosufpzYsMk5JxB/OMxee
ssX6ubLctpLPAP8UFCNreB/E2ld01AGTTJP0jBQyvjrj8/wGpvesyhKKzCgQWpN/4z/5n8+rLOoG
ycvjCWVQG9HkIFDH3CbXvbxkV2OgdbMuWoOnYb94vOB+zs2UTI3NlkFmgzk9vUQYyB2kLtjX7Qep
8Xs3AAbVr386x0h0yTQvz541Cp3L8Sa1Zzibtu/qC+lT6ULaQK2Nb1vl6MoNjylqlvlf8ndDoZXC
O0l1SIVYynf3fp4Hl3IMXPIrAyc6unSv8gGeCSJW7Sl29VBlEo5EhlFfRLagBErVxdnn9Ccu1Mf2
fdZth8EI+LLNco7Ji9qv7MQk60GtP7AXzbNMzr6RWxUpLspoQPZf1rloj39hEksnt9w7JLMc2gZ3
vEAHZuiGcurmBmZb6YtNyh2q2UTqS403OVzx1TW6h/yhEVDVUmXCIIzhv4WHfZP43AcRHNAkPG6s
zuf2fDw+URslTD7f3kePlV9F5mi9V01seW4aGewFZBSTk8+jOHz/oaZMJZ4ZuDYwqL8ZG1ZBGp+A
twitWNsSLAzksJ8PW133kUik9I0P/McddIRurlxlzh+rDAnkHVL1CB+oS6Wiy6wSChZZgxiRABBi
ZnwNYIqp/jMgR0F7Wu+9nSWBrCR89kXe5rgyEri97e9sSw2QgK4NHsTikwPhAPyVtQhAKgaMVDmT
tiImTuT1HkiNPcEDEWI+r9NX0qATcXWvw4R38OIlvWkxFzqw2yE6bYrXh3NVegYXJjel/TNyyBIR
qPDuF3OIn81v3lhWY/LU0Cy5SMF/4/lBqa0ayXGlnLNaEDTTGmO1r6fnBX6xMA/xXvsQ9qWBR8TD
JAGSXu7WYH/nlnhTLaqCz+KKIC/GVSOfql0JFsP11zVROo60DOl6IwKWSYIUHrEplFEMt+B2ccGN
tTP9BCW/6SpfCuxlwcnEnzK/gGsQ1sjHyRTRiUGBfTaB0WogoVWV+ASzaiWdOqhBrBxC3bm0+hrr
7k361+mIIGXwfd1cZduDm6tJyTdJzeJq61WeEaDtzJmB8UKaKJNDsi4Hii62QgwOMt6s/vEfbhtz
ZzBWVqWQDHYqsyj7Pzb6oeM8PaALw2FklVfQij9u98Wb/MqGK2P24LXrzI/47ntdxgkr5v2rkNbT
OAFjtL9uA6ZitjHzqwG0cQIPiuVrbllon6UzrIlGRBMjhbArQt3Oc1dcCM3NDFI5k49HCcUFXlOy
VOW5Ynbc0qAgqQJ/v8/aDCzbcr8CFrUTPK3zyD6gRcHnWiU6mHHtiHt1W+vr1YJRlfdBH0VcG31f
gmPMfHe3QM5FPlUPEynyVmq/OEMsrv61L5MzvM4Y31M+4V/MgC/Z8IlZ+ZRCzhGZnP7DdB673vM1
tCUaxuiTzp0SV/cydfKy95n33YStoGe7jsBCKPk2M9M75AYIo2hXEt+QkTxgcH4oHdojNPd4+VnY
46BkzZIQPvC+Tex1Bt1+gq+HVd87NXnb/RY8dWcmKPSvtkV1MvUee9kwWrBAcCwy9873WL+gLZpb
S41JZAHo/IbtWxiQXKpukk0cUvoaa1MBU2HHSYfrzDRP6cqc6TQiHJ1YtNvX0UnL8MOjBfJ3uwn2
750PSkgrdM2JjJE16Q/KMHCaJq75hZSnugP1FyDrecDmwiv4Wwnz1mHWsh9NL+uAzv5TubsIzUlu
h+H+4ytQCWIko9Xp9sTPRl+kqliSMTgKHwwWuIZChq2HIh4LG2WKk6Xy7Hoajw3RcyC+IhiwaM1f
swQHgdK/lKU7As5+i+FUltU+JivhmdLVVIQNIInC++5lVr81VeSwRbM2apRVN/wpqk+h4Z7Ps/XH
oeNMOQdHHZAVuTCWJkOiwf6NMU+7wZZKujk0RTXKge8WyE7x5O03gOu+lxHC3SBFuRn+9O5qCvCX
DZZw3DjSG9+nfaAnUxWcvlK0otK2803lqNxNLk1ojvrxtDnGmN/9laQ40dvqRBJ22EtE6lHz4nc5
LnIsSJdZzGPi5oYJczwiOw+NEKuscMJ6xDBPX0g32wfMiXpuX2friFIZj/FsOs5/0Z6kNkISYkG0
qTrjMXtvtUvlHgPAI/H4BYVlr5383OMyG2i+coBhKCt/q4iNbnhr3Qk/5YvPcNHrncu7e6eTzmX3
rw9SStotDI36guUSrgaEphfxTodVxcZ48sLLeL8oFqBfcjl/Uk/vgNreKR64bBOgHV0+B0gSsnBM
XBHb2VKFW/uPKIC2gv3ngv/pR8BTpcK5cqX1rAF2D3XIxnaY3hfFHCy7oBKiph/Ad8GGFFj5MO/G
x0KZWoh8Ti24zZsswoya3smdn0Avdz/Kf5zAuaCmBy85Taf+XaE1khNP0cwds0z9yL4O1MksNsqE
yyjlDcOchYmTJFJmJJ02kAWImww3n2P893qnU3EeJWF71nYAo91YtLPNoRcr/3zt1PIvJu1QgWm7
R4QNaBYoAWejrsc2WwAyyrMnHXj+Kc2WsDvdAgevDIpRdZ0aXIMJK9nXHu4sHT3ujrCHzq4UxH1D
heIoXcjHYoGQJl5sBWfMbIwHBXkYQtTYjuTqhIB5SWSws9hCC/7oCwYD2LEvvYbWLEBvy7QhNwDb
hG2CY29oDUwXUb1SC7y/E80czcS/9V2hYWZD4WHDYajTahw58NnZo3sbUeyPA3gzNyIpz5W52S7v
ewtaHNRnJ7AEBhniWo/8CpYP9Ze06IbGUh3bx2R7YbdGccMLnKjc1pM98ivFDZfmCWqsoJEudqQw
0Oz1c+l4/BNkcb/vq/v1SjjLsHZ5v5tViWGJn3lKf/IwrfXNMWfXsXuZv1l4TRdwBqKsPcqCWR4J
D/Q2Ouf3BB/PWVpnDddZhdt1ZvzAUzGl0w1CaTjPXBNKrIHVIODed4LQlY8/IBtGZQcg/R71jUQz
k+E2nXiMAzMavOtd+xaVOgOgXakbaDJnvMMqSd0i5L+iYuaTMrTjsRbM8h2c6HQ8p2fR9iCMZjl7
X6DGaYGE7ktn6ZpY2n5KaP0eLAzVOA4KQLVkUSNQCcPkAphm/ODVB/UJIO8hHJ0sWe3J0beoV2Fp
9z5PqTWMhUTVG14i/5rqZ9z4R39Kycpvo8wxunSkvnD27LvMgq04S2ZasNuxthjBiUKO+5SryVYR
+oNyeWFWn6Z0nzi3urWrBx5fFWwiiLZ0VJdMAPgAjJqBLG1qaAdviQzKOaE/Aph3qTSoBMSZLcbi
VkuhYIl6UpqOmV7pv5tsrR3BoT0uk1OgY0b4NZmTi58YM12/UMeSAOmEBTJwTMZGUS6Hg1pwBnby
eXb8q+KILuDkZWasLlTqoT1/URP4WlFyE0AUJlusPr4X6NJFQKCnthxaGLQH0W7UgiTtGeyBULCL
6qk28fjzykyTPf/OhIRMvu7JSIsHfglUC7kO1V8EuyYmayrI31bvIGqgFb7h6eUomGuqUDdcsr/0
MZWvV2Uqz2CJNrABurW8CIXn2jJNlv0BFNNBlYPK0Ou5lHH+s0MbyElvbjC9KeYsi5m1q7PjeJbq
itH/6orU1rTdTYUzNIBX+geyuTU2/Tdn58h8gHVW6EkYhUMYrEr13htj4LTsLYh5g5GnDodDJ9FA
inUPWODfmw3h2lcfksBsLFAXpXIdUZPFGYZFfWLL9iQUR+tB/ey3vYgavDlbhA175uPJLu+4ghA/
c1g52cN8X7Fr60LL4+pVl2Z19L4clhMolQ2oGWhTJDzPZ7gh+Mtq8GObVkleofXGXuiABVuztxOP
OjtzpnPK0F2EVg/P14qi75WhyDdAlHfya9Wc7g53U2/qcdyQR3RO7w2HAbprZx1oPM8QstJS5OCl
XLCPiJTC+y9o1S5coQHTukfVO8rQ9PQ8zUd/uCfouyU17P3YKw2pQppKeLt1VG3Et9vAmrNmehbV
VR8Rbzg8q5dJyfUaBtfUx4Saxh5mSxPLyR/+P2R+q/KZiZa2awRWrlsv/NtLTOKgrPu+sYhQwDHe
iTa1CHx038Zc1N403NrUVBZwscjVCVhe2SpQODEsbFhpRd9lQ6q51oVaASHPr+Zf7FxbQ1YrYI4z
zQocBS+gZeDoI0gr6OoTw8TJNi4dUiry6hB7kAQNExVbcNDDbdxx7QxfqlNYtYfEcBCJMIP/Scl/
neDoqU2vHcMM+2/t4HkjB81P/OcdmdK5W42uigWOBddRpWR9pfmIXB4c/tmyrpgFFFBbEfU82SW8
6zAeuyhS7uiodft3THfpg7djZ7WFB1t7alBJt34ruS8gSHvyIjykvpkFD77YXbVUm1RqsYAhZjC8
Kj1X5G5x4Cmnlwyem0AfQ90jGkj/yq8qLKKBjMBJiNPHtBYE3OGnIigjo5s/ycbbBG5Ygonp8mCd
iaFukGx9Szdt5pDVYbFRQZYFU4dxM3R79vUwl6lwhtDhTJDTV2yd+USjDPG8rKlxISRNjBmB4h1Z
D9Hh8zg8lup2k0AIO0eXx8jmNAFxHm9NbD+X4kQKv2bwQD3YUF5RdekhbssYV43iDpPuDIBkPlzW
6FPOfif2J5wR56rk1EcaJuQTpRu9vlvr2J6ucLpeaEKXsN96QyKjyqEhdd3en4F3Ru/3+f2pHxdX
h2nYSyf08yo+cdqvpDnHvTxwcra3mnKCUzOA2iXW2CBCm5gEz5qKJXZoWB/F2PALlmGPiWNVY0T7
8LtDB8Vcd7y4uIqneDHP21YtGsE7rCLhq6xjcbjGuetiFvhX3UALTOyh64uKvtel6DYHUUzhFYrv
29Z4pBQuOB1u+ugRfWLq6zBf6gdh0Gkx21fXIAef0/0eVYw2oVWtJEr81GMq8Sq7BVOUOOo2wGvB
rUdDW8X0vZAh5OJAJnatsF3WYYrIpFaMWQOuiyjQDhqnOuupAh3OrFGbab29AFPWmZSVLg+VFCv9
azB6k3+/uzldUfGFlu2gy6TDUhRnLk6H5Ot3ezYhBc9qgJ2q/ZLJoNodbmsKIxd6wRhG1t+EMnk/
844EdUlNGI26ww8OhqWT+Avgf80BVWwtXEgjfFoJzfY0rwaJXmbvOoOg0upmax8cQ5eAyUEcoMQp
sETuWqlu1xHqO7zB9EI8xh0AZm8qcmbT8UXhIGV/HZmK0A0vi27rNA5iNcJDJ9fYVLmCGBfCHc0g
wFDGwGwV1S80pZcV4rV47hFc5SkaSNqDf+wemrHJUxBtET0nL1E1sy7cOQTBYVpOLDm73mheYoSX
bQe9iE9HDOC7309clSGig9bwPuo5dYv8b3jzUBgPg2YUiUfvBvnbwk3ZDmNBmlF03KbHf9IDZwwh
Y0B3SdBT6b6c/9lChWwC6zW2RmnbhJNJMoacJKNERT9fhVpHrCG6N5tRyY4S9OxisoP6U+97hb9r
PPhf5kBD1zvWQAJ83zfolnQ56P/IS2ZXiFZCWHpFlN46TdRXlTIpCqhfggYk3LoH74YDF17FsyND
y2VfNcjxrD14R1A2H27W16i1Kgf4Q14GaHpJ3fnBP0kxp7WT7fTr++WtuubrqZ6NFnyYEAptkyLj
UupXiQ4ZgcujqQOaJOiT9Xt5VAqKduAOjhyXQf+bjCt8gSfc283lSLUtlA1c4sJN6XLOQnf7fVad
VJvgoxWcSvaqjiLNdvpHd1JdmOZ5Z3i5+3F/evZ1x/0ka1sXkabDknBYLuXbVMeceXFMtXo4bXXG
uzPqNv3+AeAuU6ECUaKMUkiQh+D7gzFwiuRUARNwFgMbAGyBaIMGOY5jaoKlhq/aNuF4hGiJaxL2
vpymHQqQ3XdB74wJNrDPQRDUEZXJFhSaOHRKjHmf/HBjFNQlMoDwWyuysUF3WrumSFOdxnj9FtvX
+Sd82ErWCIllR2FYuXViUlqZF33e0iEn9d3046Lz9vg8HklKWGhlGWO4+qwZpMZrN6vg7K31A4+a
YlNOgrv4B6Kp+vD1FBsNnoMjxTAZxRH1K6bXwJWmlxLI2gHnPJh7q1aTb8O+qC3iwVsSsbIk9YvY
WxRC336bNkJBRwWJ7DYHy7Z+3287Z9QnPqbpzWGo2oCC+JbJflfjXBZrrqWcrojR2d6kGYGfH7QF
j42l9BgnXxr5ObMvR9XcdiljJwKoTx00Un77xMQduRXQPU3FFHhYap5deJMOpBL6JXGGpPGwmDRg
xoO0YiSkMzLnbCDcKeoUONGeUszAWajzfoeK6EHyoujRqaHJuSExACUT2mBMDB0LqNPKLZkP8tS3
kfsWkx3gIF2yrBN2qpxwlq5Lg56YbK9p+3MA5Evf4wIPFeY2PBBdzmAowqbb+7XHukZA1K9smhnL
BQxLaaxQwAoe4QqNzeIB6u+vZKLob0eNOhq2sG9LDp9ewfO8lI4xptcJUigWLwedW38yGtinw0wN
VHizY8vYA+MU8rg8MjDSJkMsCgQw6tfBSOpBG3lkkcN1gVPEjiWcDYHslkHCFfrCWNIU8Hgjvy7n
lDcHoQWU+kroB5KBCV1s7odCe/YcJBrghc622Yz7sY/254Ea9DFH1bSqrUMgwUGoM0Bj2086O5iN
Flcl4Iinvz0N0KotLbmFLri3G5NH5y9+77gszBxNacOWagwb7Fau7DKpZPmzazjnKAtTCFmJkd+1
irYA+3gjkqw9l3TEs2xkUZ6Ugg5eexH6K3DelMRyOy+9zh7A7ur7ZTl6+imujbBLkmIGeKenivVg
3d6138MEcsQ4dWXZHusY4CEvXJ616B2VDBzz3vIR1Jd/nOSLm56RV9E0hS+2HEOS5Hyv9AaHZfKD
iPxhD5axb5vI4ktwx2er8+GaRO/hYOyr2nyVf6Mi7mSzp+7M3hA65utocBuLvtKt+vSskNFAmE7+
oYT3e18a2EOT+6vmuB+tiSr8/U/ChEP/DuttvbNQ/nAG1MibBVNBZ3OWqiOtSBrmTvZiRKFUojfx
Ha4MYMwjQaO2F3YPKFTox1oQSdNYMNYoZ359CunGc4Ardd97YO9vD7fhMvBj7K2iuG/lWuSDcg4B
z6cplRPOXno7Mx097vaKyqLnGKH5fONKsZIrI2Zboe0XsNB3Vd7GM3FVq6CoS1QFhjZPGcyAciOk
nWo4fO//HN8EMJSpd8NFc5/QyxE8e5UfDDdi6AMUGzi2m/urqNJrOoQVb7/DGnNNiHxRvXZv0R4Y
Uino0/CqSQ50XLuyDpxRuyH05CUgT54mMZuuDeQA9l7FBS2dnVfzmIF0yCY6RHT2rGr7tdAPfYmD
35RZbLxBTRkPdjqi/CXNtcslIUamyzUbh7w9HBoMryAkaAFavf3knaX/ibFWrufsfbOGUgDKCydD
dvovG0HkE9vdgLvQUavGShDPswiMt7wje+SRKsAPCMod0Q+IWSdATC+2LBiGB4oZ+GrP9bSTzOAI
4o6iaLc10dv+RK1veCiFlvRM28Z6G04HjRsbeb9JJ4HCm3GzaSpbo5FrTLReDajiGHIDGRnuu7Mx
ieWhkSZgWg83mzV8G1rt16ewxNjY3XPKtAOusYCD1bheA1C2Ah8WRRiyNXxE0WR64iifVjFTg+2t
dduitmw0YNs6TioZGU8cz/smmHB3o+8Y/G3B4Dotug+44aZl3Bp0RLVVFTM/c6dUBLp+1krt2gRP
OXcWpjr0iczBmdG6NyTXOrCgkRgTMub8ptQG6V063M2VVxqTYxdz2dwIHpHjOgKQjLmwymrRIihK
rafF2IlpnoxWDIRVktvApYqEe5vxdt+gDiv0u7VNQ2belXY9AOX+1YEBRzbACOakbs9BfLV1nGmp
Mp/m8xIfo3Y3gQsbw4GJHxm1Ga9nzo5k1KQQONcaLJG1WZIiU7Fz/H3P7vJLjiY+ACtzYmUoKJc5
cEcYZoGlNd2NTTUIxzvRaDABw9Q/lCgrEyYxPkCzeF5hKmnU2ffq7KyYxh53bROil30HEFkT05sf
7UmnXJWXZjsBVL06Ajy6SHWKaFkMOyqB6l5BO0fqcHM6AHxHsEHpEJ+9iAnGZ57UIxJ8+v2webIs
OnbIJYmuUbcjXA+/Frie7EYbW0j/Fvni4W9QLaPmWZ+qwoH+eJ2d2lx4ipY2nixmBwgL00SWDJcL
/whCzoa8KiYugKre7e0KR33lBEutfnJrj1iSk6MhyACTnrUCQSvCUKLoGIWVOUBJac80KTzJQMty
v1F7/aa9JpV2bIHBd9hkCqQRYIq9EQ4a3K9AinWOtRIYgJvQxoclas7ZqlDRgp6gKwK77GyfB8bq
8/xXF8LnzXB6IZ1Gr/x0mQZ9woFDyXRa0dTC1lnAUXoyNMRPFzcgzzUsCTOICR4+syjH/+PT3PtE
IvFfv5F/cpfD/SIGPVA0Gu9AT5Y/RC1ucO9CByjroM6toN2M5tgvfRx5SUpxXdmKNArOUhZ0unKZ
MAJ4mK50kV6xxggLIv0Rbn4M904ck0Z4bjGu6s4te7dZxpScvsBnHgFD/DC75AU9B7KB+N+Db6gZ
0l/zEAqWJ1T+Qk7Hh588KS8S1DdAPQU9EwAETh2nTIykTKTIKDTIQgNDBC6pJ8MxYBTrBzXGhmvD
dgXzN2T8IhkSqpquKZjRw9Tl57hWdToU4fbuFXhDUfaLYHG4FYDQi579RP5ouxZxewqCpQRjfjVu
VQWNMdnFeJh8l8IkS6h55VYQ1Zp4NSKtcj8FRChEMN7GDYB0OJkNp3HAX4tltNINDmFXlY0MKoaE
rY1GLOPhvpeVkeci+dNhXdvSjObMZ5xavQ+PX5/VDRMwE3HOubt2EOfFl0zYWbHo5t7vCLmb1rdX
71beXd/TC8hOBxyXo1sSAa7t4p2Fz8bkut/MY0Ai26us0YiG2WwcyAHoDCYYQbcMsGPerUVJZsct
dnMUm/8iQFku/cs7zSkdD5TTNFm9fO/dkpSgYYaG++bQokNrwSUuBb91g+Ib7tb0HOAkgAmOaMuT
rw+3rj+RD3iZNrPrAdPc8kQtv4w48REj9GSQyuwdit0gGBBTObMoYIExcRVm/ONma+1L/5wrFqGw
+FtS9XxwBzNcAd+/2Mtq9Qv2MlWRokHtCDDWYi4bxLaHPgfxSMifnQtreXMcG+5DSweQAAv3fHBX
0zLwQvcBlQdGVIxkaHXDbjIAzYoe+B4va0YJZxefbhZShJHnJnHNn2mU3zhlW1kpFIu9n3MnbpBv
lvu0OzNC8BRp6GKDYbHFSaW151zgSUqpszbnKs1y6Ck+3g1KagbMkWO8rUaahg9MP2Bwl+y57RI/
vIKYOLLi1+GT+STrnZjfLSLCvnXmBiS0vYcQeiEAKOcs5+tJizc7ZGN4RTNyfOaxkzFyJ+GIu3pH
+TysCgRYl9bQMGVEW8sDxHFhZ4D2HczDGYAGcvOboZZxXzKMMu3Ubalc9rlOjfDHopBkFrW/pYzd
10KjUy3y+OJteskvINsSTt4a/bAyvr7Aq26YIahBUR43be3O4NIcmZkd5P2N3RmVMRWa4GkatrEc
AjSgN/6pjSsWlP/5pFQOLdQMlDVYYbAb0mr+HZx4lDODGrWkGUJ1tMoouuRwPbwrmDhCfQ8EwgsT
wLrdI8oHLYaJiZSxzPgVY0wpkYx4sz15VO5BmRWEl67cm2p6LHbbLrVoW9gvg3CQ+RqFMm10UQ/E
M46ohbuLrxr1KHvbEtW/BXSDtdDK8+Hm49rk1Qz9IlbTjFwtUKRtFom50vfh/0OvBWcOy0cEBHTj
RHjhJcaEsj1SMUx8mYMyZlNhNpu/P4gEOVEdPegiSa/jZcYiGZvVAbFNGnhQkJ/G1zHtEEnp9j83
EJh6uvFVM4F7AbacgaAxrEW3KUCfu70C3QFwAoheDRGulBcxq+Wj6wNeThjzfJuMJy8jHj+xjlYp
JkSt0No/6yOE1XhqcZdDBuw4E9fECpaTQBF9w5kwF+j0j2OOWh/3HThg3IZCMwcsJNg72YnXMjty
hg6odQ7u/ojiv4B7K2ynoqh8ih1Wr9ix0v3BsiBUW8lNHkMlV8v5+LsznvFVU81Qo4JtVqK5WBpW
shpSrZjaTSX1zKHsb1axnrG7rvVo31yusI1Ma6gzNVKmzstGPqsgSl32UM6/ASk0j6dZaD4yShEl
l8zsE8LRb8vEniV8e6jAvZv1Q5U9vqwRw+2phXt8N+paxrNY4VknCaYMhsMOy4aDDfRi2T+J6gnV
SZGs8lGx/ET+fh+liq2iisfDOgqB8JKCpxSM2Vebe10vaX5aCwPRGGHRk6StPFeqcxlvxoUWwtQa
0aJYF4tKFX+KwOMiPu2M88N4HfMbNpI7svnXrbxWgKfqlVFx34Yo7e2bpgxNZJg0o2zedKk3cZKH
ih8TDUTC7uAspvQnmtBAU5v9aD/t5Nh2ec9ZmyGGqEmb8ezpIxJHS+L9LEQDzJc6ql/6h7E1jjzF
aytuXjDiq9vEuAiR34OIUOdX9DkAkBdvVM9e5rDnhDTNLIKoIf0BmQVonubcyu2yoDruZ1h2c9Wq
QnsUSOXN0sxnkBjU/MvoLntjWktEPn9KNbX8UwfvRwuV8fNuT2WGdSfYAYpfqAEKEntIiXk5UsOC
g4PpKh3MnnDtkP6zSgXRUeRc3d+XdHiJZq7IJsRAeNRs9qt6/cN7xBftvEyyfZdc5PBCyAifEsC1
wq01o8WsnIkqgEc6WDimbNmpgVY1los9d21F+wULf5jnxQtPSO3GTVnZYRNWLu2iMwz5jxIB88zl
sUuaGFbD0oidTJ3GsOtBx1IvFZXou3oaAliyerUc4mANZdMINbO2Sy9A4hoB3ZhNhaUO10r7ni2z
3jjhflpCWGXAn4k8eRpvhrO5XcPvrgaRtw4FjbpaVHElMJzWknVURdz/7cr6yJ8btBB/rl7xurL/
blpeS23U2X+Y+OXXj3MrgisVhodAAcrqhDXeqGbnM6GjMq/41fIhERgYPZVu4GXYIHaNH/Gya0e6
p4utbbf1SYZKQIgAKMNyCyQIoD0ednELvUp6Ym+8AwdU2oF4GjvKuRZOIO5L2r/4AwlhtJWdZd6U
vWXvsxhkZCaxdgUwf3MXYZcFulaE4oYBMBieXml00qaVgwkrBGjnyZOWLX/dnzLWKev5559btGDL
vPFTmw/qA+32zOxxwSZ2CIsKwaCF0hjfTzR1SFBfV84r8xkTprP8fRiTkZ7RKgXB3hwXovgKCy3J
zY48gcS8+Nf8iMja+QHPP4W/nvVg/q1KBHMk+1mcfT/LwfGjn/LdUQ8+bv8O2vl8brg9xnmQ80Ol
4MlcIpcYSh+P/vM3NE2pXk0OPpPAvJXdjKCq9wVWzH7edc7eRSu6XRciLB3ubodeYgt0+eWZukCq
jMavCgCGBpWrYdcl1l1zW/dwNsRqTnUifs4Qo+g6Ga9dyaaah80cll+LqwedVaWPls8xM84MOyOu
kyIj8rly1jKGg26lWyjhzNDeIl42KGmKFkuz3OKO4CSYmmY7b2KmVSP9j+CEfLYIS0WsLkWm8tKA
Qmp/1Pq7xzCaPPmSZxXLNq0o1NwtaqoXaFLBuCugzPLhdGVimRk2Bi3cyIMDgp7pEdhzw/aQQmhS
BxqapyXgm4hSX/e4RncGbkAtm/VNh+YIR7fY/eob5MPAg8iHhvOyGoerwmNaInsZbs9px8YMrpH7
rZoPMZTIeY5limpGzHVqNAlgY+LR2RaNM4uNnwxUwgHmga60buJV4iq1BFtc9oJ7ctdj+HvqnB2g
xyc6FXXtH49kITZpaLdoyCFalR/XVM4f0w2qaDY5C4TCeRpZ4biqwx8LafTwu7hotatVpvA2TZyi
tQrhT2/MKDns049/aST/fzPCXh+6eOtbXYe4CNLSYclWNgf8WCzkHjmNeRGBexbnmBp726XZjIIk
am/6woRjX9RhL4eGaFxhsIdz7idbP9m5Y2p2BKGZuxahzNBMVi/tTIAKzmu9BnX65cJIMlTzsc5O
6fpVpXdJWtbyykzwyP428Y7T+Gs2yKqB6HVubYNoACyHRHVYB99Hathz8vM2DOjGrSiuQMMvip7a
bclTJl79VJ853lzkV8FpS/7ahklrMBLFsnlNq3qz/3HYgGogifBlqHEV4m/yJk8oDKNI1ekZxYu5
QXLvMHJt7QSsv3XYw/ISEzDJokIrxhOuTqHdBhBNvHuwnE+iK0NjvPdfuYDElmRO4pT9KOuBVlu2
Iw2IUD5thtxLl70qDEw5VPqTvPODPhuOkMBT1WXdkdwXTZWmhbxhcPcNK/iy4kN/ucsPSVkgnRr8
c3EEtDz/wXj2HHLLSjrwFbQQAwTL2w1ud26XXuDaGIENKwj4CKpWOJUel2i6HR9C7QALg0xhKds3
bAkacKff5uTR3FjF/l+alTKaWYnfmpGma2QNYNxAhY+ZmBFj+5fPmZ1wSLM1M/Ji8g4e/2JmeVPP
UAHV7YkZpUm/Q796emndRgownyJGFh1S4RfODvugoL89JDtHBzmhrSLspK4rBuPRo7B0v9Jr/hoO
dEpkC+tBDpQibRFszrhEATRE9oCi0OzCwjUN4U/GLCxLP7yQEzc5Ty7MHJXEa76XPdYHlDzTouxz
5mZ4Ezu8/iyFIV1d08jzd+nKlCbiUCWxm099dDzTxvl8KmBQlPyoQVq6xDStlNt77dpJ5bHQIHhg
Zji5Xu3ujCDYDV6qJQCUKFic4VA6G5vFmHO1YieBvPypgnZAPlQDYl+UCl2fkzkbACQudAPwkAb7
J66QakVbnIZgHYs+ISyyrjF3riv1UbMWX4kRg0D+6/t/pj1psJH9UaTW99fIEPq7HYawMLz+JDq3
zTeKLv828Z76dvdqHQQ0RAar5l8BPXnK/xOuj8Y+7G7NXDh+LRaqGlP5miRdbGU+iSwe0HtpY5/s
dqPO1AJSnF8oMYgLWULgYONz3xj3HELQaBLxGGyQWs76f73/oh38QTfBYZGKhnef3PxmmSio20tE
XiFj+mhm11vGLXGq5Vsts32flyTexFhEeQMNPXMLHRbT9ghIwOtRV0Eq464B4BUfli5zKNP2yagh
6PdHeU9dsUht8Fcz2duUGnhCwYtk+47gE6s8bSkiJkzqCP/9RteULSYel4N1oX74iB2nShEDwF2T
nr1wy6Q4Ez+ykVGqZRPi8/pmUFuKkNDFFbLPGvkt+MxQAWUDugC3dhRsrRH+CQNQrN1SRbMvoPsN
rxc5KmJfvJLDZQkU5NPkoDn2lrCdBhaIaR51/Jo6UBFGkuguELYCPpLrufgWPfqgjmRC602FtX5K
aSguHBwGpYbraRkZPl2mmA9UmeAv3i2jqbrVedeEFbKU40MakXIEz1mZWQVlp3QR+98ML8HLDGr6
mN/cUP4kB1lXLjq+foxoZ1EdVMWzs4A3Oyn15f9QcHPymYbjMVAmNKs4wN0QWKrffonSGyWJmQFX
jPJ5ys6AFD5dG3FNN3J1DUNNx5hhI6Qxbr859Iq9ITYtshjsTowaPkbJ0RSUPTT//u8vs4pZPVHJ
qDNYNSNwzNBVFXGEPKWGhJap/cWrW0fPup+Oo2H38vdvLhnHNTXbAPQrwd1WcDAabEXmpx5T9v0t
119J8Ax/hJMih+aqoQRay4kS13vs4WIb6+mH/WWGzuuESbrpDbNOX3MjAh4rf6wQhWntKScZpnCL
p8ZNgOfNkhziHlzNRaZcEmjyB+yI8gB00PbXZw7r8WMyJ2bgrWxQqriGoEWT6XTkworCCiW+E7jA
obLhRvovC5rAk4LGYBglBlz7HrvCQJ+wrpCCmECwIpJxG19RW1T6gUHwzzdqq4bjrtDUwRSHH04X
0gb+RuU/7LMWNQhMhaI+H8aA+Gr6w5AcTlahh/yKgSMTSqRrvnCItJ09VfjfCp7j4iEmDOFZOL9P
Uvd0V1TX55MjW8xh+JgOWNQs58vXHlyYYt5kn/VlYrDULKb4bcgnwkjtj48g8veYhd11bku3LMrR
/rPMmYTW4tWeHO9r0qGbz0kyuXmKuMnepoKnCqRtMEg2qQ3B7+25IzPRHTTZzt48HG3mg7WqMWTv
cKWJOyQw9Mv9JOto79SS5oalcxWmMv4kXUQZPGk8Z2ET2Rlct7t5g38xnMxo+UpK/2N0VXf/49mf
QdwxpUGSNdlTg3RO4Me8OfHh2LuOweIGICG48wy/+cHaoD03dspS0BHZ6CFIhOBKWbfEvMYwhMsA
CcCkReXg5TnlsjhvUL0jI5Dg17y9aLoR6cEtY9TwCHqelAH9soDzkGX8LlZ9Bsebe2pMdYf/Kpgi
/7fSetlTkmDN+XTZeLx+LNIboQdnunNFtJakiPzIpIVnrKiy4htrBNlOK/zRXgJnhRdTcdNPShYw
E7HKC7ULn+JZiS9HYv/OP1/S/4P1ohLpUtyiUkaClA93T6TxeLgOG7NGAR/L0zkZjiEFcnu6Xz5I
blpFcJrpoDNQ15upcyP25Numz888M54Nryg58oC16Q3hrV9LJBtMnSUX4mm6wTFxXwUU0HS23wZp
PuU/4sy42oMLqz3N49ENXTE/zxV1e8iDstIw18XVVrHlLDo5wRfW5uiE2DGF9JKhQWyEKMtyOxaI
Rc+rWdoAZA43x38VaAS4XKpFvaWhVelAJwxa8b+Y9SplKHps0grJ9orsUkmlp763hbvg1mBRIdk0
BP/9WQRGd/sD2IDrXoLPx55AU9gaf44cZZs+w/XH3zAcUN0VeB7QiouXOVl3OzXiiiJDhLRzhMfV
sNCOJU0UpYndJKUEaaQZtRBSREylMgLDfdZPmv7WqZHJ67uHPEn3XdQbEmGcWUKQBLlzII2Sd7+T
B+WBxy3lhNXztLlFqx0wwMEgZtidKVeEIVE1iM4EcWm2Sp/wKyj1vuAA4Llz+WF28C4D59M1uTQr
0bostn9sAmyNUj9WDqJcW1ClBcpFXqIkDNZdGelH9GAzFliQ1hETyNJ0pKUQaHegvo6+nYSfJrLo
XTQ/OPSAjwkXkuTFoqtTY5aznBTVo6eGY5vjK77vHTBPcW2XZCoZ6mPfgB0NQKIClzQbt2i+Pg5o
l4zJZXheD3mRu2hUrdsc3Gi0z4wj80GeFMx2hrxO4heh0PWqD+faXe00Ar0py+p8y7sBiNZWDgqG
TFlqnTvPFa9BSw1C+B9vGiZdFvMA5Zyhivyd9a52abrEpwkwPXLvbB34amKfX7aZfrLEu0MaOAo4
GH0xLg6AFnNVkEN/oAqV+CJvY/1MtlmR0aO9CWh6Er22WCLbx15otCszXa+xbULVwC6EmEgbxrea
9li4n+9u+BhW77hzIpkVK1u8X1LH8PuG0Bir5LBYYdH5o6udfibt/ID2MdQiuW58hWmr7pXXMH8X
oB4PAqeoA8bZHRs/vreXG3TP+stA4YRMgNBfRs56n7OVl/dmtuajFpJ6q01s85VuoVZNlIhGikCW
CbfnGeGc1DNzun0WlWynZmIK7jEB2y9lVAh7pbZy6ew/FFwpi4ij4KrAiDEw1J4AzoBUebOUQf/2
qIkm9KtOb6apbPvwKMjXWuaG4Q1TXu0jr3uUCdcVqOcJK7BsVxPGGJp0lhPlMwBYDHO4d/wdYehm
qts0KXLrrGJee/n39rbaH7Dd8CcnLzzCpXOtf1xc7/O/dJQFNBHMOXuJ1QP8hp3MYXU4XJimGgPM
8ukVS5SrNiU94j/Ynoyw5zRCleWVkTogMlp750EGGPi2GFBYvJ9GyHF5l/SPNVa9eWfIfhBniXzE
Uk7Mpgow6QVPQ2Lb0+X66l479t4aD1eoreYEUoZhAuAQTOjIUi+mYqm9mPn5YfeG+8Uqoqyn9t1v
UTMXJunrrRBP0oA8y9PmryPtAiXl0RZgr0qdgkYyF0JM3czAB6Ghtx3rzw+dkkMLEj43E8ENkLao
V2OpP2C9MFT3PzQtVG960dzMj4A3Cj/5aqRcW60Y0A24uHbq5ivuPokSJb1TljqcPSoPlDe1xZN6
XxDjk3QJfrohQVaFj9TxuIjBSCZqwdAKx23RACX81KOwLcBfiODGaV5AH/JCFfABZfpXylLFxv4W
rfGwlfx6220YZjRDnSlLtSYQ8426bP8r+QxXRUStTF6NnG3DlJ9Ny0NPU68ULP+NKR3ux5srrSuR
0NarXdCcre2mvL1jxsAVHGQ1K0nN9VLs8yecY5gXhb3kVTGwoUnxhBoQ90J0umWrK3g/f0t34fiK
gniuenstDYH4y5BKo9Ha8B1WPqr94WuuhCI+Vrix8nH31847Rwei4dlELI+6xyLvKL/o+vzmfSUx
njbDc3Zn+TQNGDjvwrskAR9nQH6MSkEuWOsTcmSSXA+ww78ZQOYBVDvGYnCrXRwpUUiep/XUaG1z
KFDxxZAMy/BMANxIWf7RunSmT+PUOL2DmCv+ptHHiV2T0GCasnCz9cLtuRdIRsLG1qjCLZ51bTbR
WlHSo1ebCjdi0C5T8tPcHp7zvCLlgn8IfW7etqQ96YAfM9VMezwFu47rUMDbQowVD1Xn/N5G5zNW
i+ci69BtRGUHtO7vuzICoi6fURsMoyA2kWKwbiXeDgQUhavNp05hrpGeyeHW1zK9CDnGuD61107X
DcnNCSw4cNiwcYaQXyDYnws9YGD2t61fNZiN2Q3aLfTaKqNOgWw84tiDtdtx6+tgfhAeWhH69ao7
9oHHv43Chjo77LwQNFayssN7S5pDEWLZpYQBv35uYEEOemvbvZKlyVlqKAJH71gfQ0b2iGGLABHL
UnEQHL3eBjQ+30tEUtCB9YuxFTaw8HUjpWg58b4mbUgSwADrLAi2Hl4cAoDbFX9cNwJ8EWnEENS2
xseCfW3FiILnbmJk0bj36DYYOb6wOurLY9KpWurA+C5ZqPCugK8LfDcChl+QCv8L5DoKO+tu64GI
xvlqtSE34FpYFlEHN61aUnyg4PjN2owRilvvDS4w3pNW12gQP71xrBdj5+ol06J+wlz+OIEp+c1a
Ah7b5pqR1pCnFFzbA6IgI8Ud20QaXVtmv9t9yNZvb+7pMeTLUag9pKtd+rFJ32n1YcLUj1aQ23hM
+aeJNFnl+1Jj/6Q0uwwHU7pZHq9UIuYOWwgp/BU8d2jBkGDy0sluqWNCANU/fgW8ZUCL9ypm07GM
nFxMJPhdEkAQU3ukK3CC6MWydbfhnopLYgZM5IqUBho3e4f2XwozHapV67WxTSV+xQMTbdVD1xSy
LMrriLZS0fJ/lcMpCt2rZSG67VyIYfffUI5NIYL1W2hB33UMQxDOmaWcTh3AUrIgr7SOlM3GXEYd
YS0NOswu8oi72lmK7A2/ilK4zXAknscaVR7TljIfxWmd0yUjpCW8RH72zP+DmFEiqZhHf56LINLk
jD4LM+r7t0qfNDBdqJGvtrnkaoStR+IVjRNVBfUwB0zavInoE5C9J9DPV9tnLlzCVgbUeoyX3qML
S6t0pGLbUl2IoPU4D1GCKaW70p98kH3VN3S1A7AXDTuMH5GpIDpdAJpuTWBIotLQ7VZwE1Favr/E
PoudYbx0u/K0S+y4NSBSiTCL98y/aQUJ2nun/HWrBvs9vnmf5qOgnlQNnLtK9ak5k1pcgNFgRwdT
UINoEgMAepGSnfJDibob8in8Rs3xm+hmnXfpodt4iiOUi/GOr3pjUHufSx20yulAimlG5RVb1SPa
iX7uydwlJ+/8lP5/mtP/o7jeeJBnljQzWS5+jxm/NgrVDfVQE6UsC9u6FyjNdc+UlpdhmHFb30Pl
jrEtaERK3Mzb/An0QzAdUpmSqkFhDjrgaXJpMfbBfH3eS09cH08qk5FuTk/5ClSyWmIUYhkgzrhs
URCBnWBDQ5QMfrDAMHr7n1Mgw4r0ccANIAQ1rYNSQUzX6lbbW3E5ELJhz1U0PzYJcwXPJ3rSpt1A
4wkcNfAaC1pd383jB7Pdq4Wb+ZEfd3X14Bx6ZotsRujBK8jKYOMXRmbLvfHa8bJpqFcQ9LRQDh/b
NC/1ffmZteLsYtK0iOxrGZ/RIb90SmAbbVE+aoZYuIt24YBo8JAIk5tiduO7YmvnSGbeqU8ABvxf
kmDzL4z3eKfGxWQe4mWg8TkFLB1Atlz/rUtyPNlwob5fOIUf4TvjOHkRA3S7qru93fgXm+l0HY1D
4ssQHs4QaTfUTdJY/b2cHUmWgD+GbE7LF1f5Fp9ad40aJm+LsnHelIjeeRZ0uUqLu3LENT2akw8B
zCf2mtJWNEFeXs+dMwPUiQZxSpg26YKmXcM6YNR7nMTZIEs82r2WC9/ci7NoWgnLHFWPr7MD2JND
+101+D9/WnoMS2ZJ1iel5vwGdRUlES3RtkSSr0g5redhOLf5yRWo8FRaJaU/nevgUS/DDlxSVtRK
IZW3vi3XJY+FtbzHEubRYdL+olKGPUyre3gKyr3QbTbkTrv2KzQZ/qrBKPUtEbCPugy7M9HeB44L
69deGYWsxkXopU2eMwvFmKWsSAUia2sa5VNG1fkGxBxjLZjAO1ICKUpC6rQ7D+U+i46LCXu504LY
m8jdjVLNQYnwjnVvTAYsjHFE25t5cXU64P6te5iNwkOlfn5ZQyTST+mNu3NRoqoMz8wuEa1ptp6a
kZmHx19aukn0qQA7+a422L4P9M8WXi9FvvxJXXezEGqiFT2pDu3oJ76klblbTWHjuU7pXEECnpaR
19xVxnRKRTaNYochCPFbSAf9TDEJaqe3KXR82fm/xxlzwltec2ZuyBhDWCiq/KHM9tT9RpIkHTrW
ZBkUtX/KXoL+3GL2fL9aiVa0XnEnuj5kBPrqeef3/YdE+ZK26FClcCmfjtMQwU7twhUm+uvYGHgs
GX14Px55gt83i/H+W0oCb7C1SpLBQZb8Y7tAzRb3sqhK7HVqLT6HUb6Xk689Fd91coEeLrQvsRPQ
/q8PZQxlsazqE0Ei/7hh/EFtsfEBZXF8NZOIG3XB0YWuw8pYZVvzbyWlawg4MujajYCiHlG8vNl3
GdZL5x3D/pDzu0BxTtJxYTKHIplaSknqC5nh7bWuyF3WZF54HtiGiorCue+mKwVpO2vslRiwASAa
NWhZBo6IlHswgYVHdEORbOb+F0h5orICsCw8xZ9hY5F1NwYcpFwE6MpkMYTQOvYfikzp5kDH3IMX
2EEnd8zHAyCeykV2qivjKTZxHFu6WpZAni34+lhWjWbnKvxlgaPDrJDZImJs2hDmouuUl9+oCzZR
8n60kx2s6nmENwEmPwVa5ZCyraCVNmKx2m/+MJBj7IMHe8aU/Ti2vxa7yGWj+PHXiqpNwozfHL6L
Y3/TqOlTPXYfFTEuTd86zEQRXQgy7YT6wCLgPtHXMCimbOrVgMZ2GlagC/aelIf0kqeSvVlBOCTL
37+0Dda9XqT/tguva8LOWXUbDxY9XX7hfOEUHpp94+QVfNrrETJFiOWEa5/I0siNRf3Wzzx0Mwbb
rKO7ikTNbeQwSLoMgisIuXR559jevMqP+9qbjo7Xowd/hhg2cW501YEth/omyP8TLp8i9ySgBhvj
BfzysZYY9xavIoFQkV21Ix728J8NaRWXVMorTTjnC8BXtFcWruY74tjdr5lz4xo5WDcq2TmBhT7L
zS9LWGNtW54/lihmuOymY2b42YgfWbqlP0eKUI35u1kzi0oKsAnd7TntWRm1Ws1hSu0dFmgfHlt0
E9rDKj8TO5gtJsvafm/6uQTZSiBNeQ4jNWdO71MJnjxROmOop58meU0Fmhx1fssJ7VU07kAukfaq
biP7cbdyd7Qn6ethlDtyycfMxkKs8pnujKKoCy92LWtdRxbeq+MAKa12MTcSVd0oNpG8aF+EZnsV
W/CUQ00GWy5VoRa1MtGsy9DJkHPwDx4TTkxgcOCtaskHvlYJzehFvJTkzLRD+lxbkWVrdkXG8/cS
63IMOBfYuQ/MsQQ4iHy4u13PGtfunZIBFUDzYH24N9MoAYW9MKNWqdQbo73w8VhvUfsS5KwHerEU
/q/jZidCIEywezibLYioIAitgAL69W9Dhpk2MNPsaFyhfcSbZmenY0lerBN/50VIQ2q/d0iy8JJf
gpLR76OOr82gRcIlpyAXBiE1Gh4iUbdKPe3+EG4eQe/0E68MIForEFjaYOcAtkS6ejkTI9RK+tQJ
Y6Uu8mLoe2LAn7tL0aEnm2Exs/Ako0kc/fL08upEExnhnLr9lqGNb3NNFkLWSrVPVqqdXeN72oZz
9eaN53laksagMOzPBbhvoqvSJI587pPRD/xKFv4WCNFedFSAXN+Rs+eZCOsZBuktK3uIuiSiD3NM
FHVVQB/+OA4B9GKJox9hhDXOuUHLD9MXvyiIbVJhJNLfKI5XuZYeOF9zx6DPJKRoaqy+yaSzWNCd
urGDEgyAYN0NS+ppeeLb9dvKt+ASsJEojRtwPEZcUk4qqK1xKbQ1gNMvM1kwCYGjhjPPI8u5Oo/P
C7GitfcEOSOtcwOQ5R0/r7bY7CMMS68y3N9Ufy/6/Zik7m3YAxmnbU3xYQEbADxJqvU8X5OOcrWQ
IJD6v1jGiE8jImjweGMUhb9lBQYvOf02ZmLeOyDaG0FwDDE0kIn2p9jJGFqSoBtr/P8KqH4hmnX7
h9Leu8cXwgIT6QW65KHCV4Pz4/wixYSPLri7SI9bl/DnNVOVjFv/+tbBJVQbZEMi2Otb8X5c1aYa
NwHOzIWEQe/mmHdM9yXpsrAQh9eXDg15xgeqzdV+S3iCZqYupnDR2A2Cl69lT+pS1bwdYFSDhK5P
kSppaCbDgP1RF81N50FccM+eYtCtL7zCfzZ4SvVE6JHpkc7nN3yGovZ3+2WdHmOaaGzpmNw7bi2u
r6TN8UxofbDXXP/V8wuvGAHWYQMwjCoR2YLhOpEANKkXcz9WjZRLNRfp/VfpDxt8TVKgBgScfMot
VFQX1pcvS0eJwiLolHK+Y5QqNpiHEmcPEdvFRyt29quyBiYjCd9Iv4igpd9pTod1A+GCuUMlN81t
h3JPGrB1mdAdEwsCQkszqdeXE454/r49qYaxxkRrakFhSV56zw5SA+O4slMlwbryGsSJl44ken9K
cj4qrArEGoTJuXyNdPLAkWgtaWbe9t+QOa306pryhnKkDIUKpIQ5tALnEWi++NYHP9YWmjjh/yB+
bdqHC2KVCdXihiAg8KZa2x56erO7eQwkNmFU2D9c53542BDOhhgiD44UqAsHsrfNc1+MauV9eEjV
q07m8JkTstpxHKsjzbJRJHNRTj8AeZy9yyxieCRipZp6/Yua9dSK062tb2kiuTKvTA0TtCg1Bydp
hk5IYhJsIWtq7AazGmUMJfmF+pMs6iMLfRxKqmA/D1qclHcIySlf76NJPC8/YLk8vg4J2uwcK7es
T/zJ7WkBx0pVwTsjnWd0Ib9ioHYXeDie7AaYDoJzvV5bkP7HjTMpu5G+8UaLRtPoz/jWn1xZlPrp
f481vY9XWKkoM3kLz9+1CwRylGKajL64u8/OqjFN3RoSiRAiD7nfGXRd+tRXgnkkNYnmZd6ku2Yy
ONK0sBpxEQyyjREf8bwVGqGqVYdwXs48VETlT3KSh8ejEcdYXxFjxmfKR2+PZi80zKTgQH2YWIgd
rls8NIJNffw5TqY0NfbU/3wVJCz8OCgFs/1Vu0008uCCr/vIdwzpoO6LM1cyFwOrOk0RYxmmXPew
fql+tB2TAZJDvfk+K80xUaBL3r7G0okXsvte9NF98JsIqHWqWyAAGBMwwsqIUy+jbL1lvNsCR6d2
knHJ+CGzwlsgwMHAbs4FA1YCj1BzLPL1ivJNLzS6goDo8gkSqf9IuH0abKieCgmDnIXeTv3ZpTmb
fZv7nOFuEijFQXukCdNkkPv0vZpGb5HEGSV7h0gLVEQF4fWPigQGx1Mi5lsNQqYicZegu3Quqg4W
jugydMauPruzs3KalWvuvzCfy73LxyelzkMJ6aZJqJe5Owb01+mVWplouGt74v8ZD4WqdfKbZkjB
W2jPdEJhTYO6jUZIlOWoYqiP4HdBWbjkuQJgoS9jBwVHHy1UsAqbJ6oAdEREYONBqnV6CA6RzbQh
WuOIisWYFLamKXWP4lKbAPx+BGLpMNdt5R2H/epb1bgOES60V/8rftLVEeO0YnFdcqbH1wrkJeWp
VovM0KYNI2xFhdfRZWAuk3R6Zp24OUnbKqFotw0k3QLLAx8OGHag2Wvw8928z6Xc7HsE8ZbK3LGz
uuBMDaqeEngO7aAK7OkN2f5B4nxinZZInrGRXAPTz5/xXhOS1zVI9fUzUnQd4HNMix8+63qrXqFz
HZ0a4C0p7g+oUBZrH/NpmhCs3vU3X7HsMwcl8eGmzHyeJyL3G7NLwuzwIPu5NXfCar/IeDMJ5EAk
7WoCJpx2k68moLblpmo3eIE+7m3+lzHq6c/ZKqkd8m2tpyEGpLcGcchi31RjXk3cDrrHUVRs1L4P
mJnZ/ZnU++BHtaeTqsWW2FGk4Mz3gSNwQnAxhDC2IG3kWzXydDEbopA5Q9wmf+Oyv7Tz3az28bJm
PzAhKqY6oig/gwF6D0FnBuM2xSSD7H/Gy+6CYaVQb2emlkbqPIVNDdAj42yVud9PX901ur1SCHqS
touF3u0gIoF4rSai9IcfbWsb/7F9eEymdJDAxUfxX6u9BsHcVs1uUOgKRrF9ug5lB+y0g5nztL5n
uAtSbu1YIJSRnA0HcOD/I2BJOEkur7mA3eTs/jwYelWlDwxjhCm55DhKfV1oqOPxVaLh32hWWC/2
wZyWzR3pjxEDvgFvJNbw3H8T4M+8wkCCc9jAc2QLdAkhUiZ/Gb95eqzUs1nX0d/Lx5v3y9PPsHWq
CbmYTQ8VwaoEe+FEZcwpIO5jVxXHBocKFbkHHMfXXgIpkzCet+ybIBY4yLA1oaA/+29hjNjqckk8
RXFq+T4XzR19emCJLx+Rn4qLbsqnmzXPYH7R7dpah3kaP8GVRrdaP5wK4isZsuCrR5dK7wOz27D7
XG6ksU+lQL5IdOP8hEBS+MpX0b/NumWPnlZWCt5u8t8DJGHOv5EMSyu3/KHB4v0aKWhfmdjR2CEa
MdNhwPRaZtNHqL5bJqj2mygsKRUzn3ym4MdGUs0y3mLflWgiku/5DaE5z0YogG2NENNfK8lseD9s
t5akoAnF1BTu2SnanetqVcLWPHbnJNYujWPFq+i2eRki1bFC87WR9NQoDbgbOYkFrCco27Ix7pxd
gqbnAew7tiKRQdng7xZlDf4SkkopAr3maOu9p/UpEpE287ihBHFBmqLLtySrorrZP86aNo1eEYjS
s9q88roYnt0QixSS9k8laoKCSD7TsoPE3LyMOX/3f/XrPglPvPQ8eQld4MJQnMnhaI0js4AK244W
/tm8BK7E94+mrGUzfsTzf1Dy78Kb65OddeBxZ46gGwO+EhgiPH3KRXmHRUKe45sgJI+2gjTx1fKU
5rmkrHTqhYs3EHKduMkRU5MOUp4ZoJ9rpZg9bFzftnuYiQfBK/d25tlgp2KXE+WV/qJGAi3qBphW
+MqOg93z5Y4kqGbNPReuHyQGc3fcbv9Q7IfRaY2cQPdSg2IdjN4ETBjd2imy1K6DCPw9k0+StOio
4fkaAiEWRUxAiWN2NXXnmHOvxtUcfMhki9L4djhBmjmiJxoyhbkZAcbJGDVBZOU5zbrtWrhhuX+U
hfnWyRxMng3YBqSD4mEAlcOJw/ZJ6KU9+Lj2zqjEn9bleT34BRFz/GvfSXm7sSTc4Y0Clgd3k6nc
iiIW/3QPxLKBDZ5LBY6iQqo4nVaJ3BbvUfzbumnot0E4wESKnb6hZSipIgCXts82G78VY1xFLR0S
dzd5L0HTlU6L5jKKITYyEa8L3PBUHW+igSN2MQu+19EUSTgFgjv/HH3Hlplf3ewEYkrekVrq+9g7
LMn5wjcokRSVueCHXCeTM7ixtC1fAhYcPoBwPla/knN9+mkXcmeh2DRYhfAvzZb4pbnCott8cSrs
UKd7VaKx7qtuVJh82fQT7VovsbYkZzrFpHT4McE5XHvqaQWu8QeDNGLZxeVQYO1yW/o85CImVP+L
lPGT8jNYOn8q/ryuNOrEFc8ZHUxeWjJ9W/MhfUWYbS8NsWpvqJqYkB7g4hK9d1xV0fVxeNBUIA9c
HFaDyBDJrPdMB3rr9e6HvY4rfsNBYvBkhrfdWihwdkdKaJ5RmOpyOUDX3ieZNed2B2NFPDWCmTm9
IKY1fxaBz2acpggufWjAjPiTzVw0YXPcnf1pdp4xuF/yMFk2uKqKaAgeDdxfr0fO0PpBbluzdR87
HNp4tyT6iSo9UCQHc4EB9QGT2mYvvVnJiCt34KlhhQmi/3FGxT2vGh8beNCL4cMwRw55I13Ykt1O
TgRBCBZyT2lJtvQfc8VTObKs2x3OOYoFB1wu0PwyGeNO6HJ5lIVfawto2vbyWWmt8woTKXps/kIN
Oh4QeJCpgondES7Mig+zaHi/8GaDwYGrLOPmZP7n2nkHIVx31AHrkzV9h4BYekga2g2PTcO1fl8M
CYPEQb2qZqI/o7c6TW435QIhrKaZzAs43I0dH29K+87bDbO18uHN4MlREw9kvLcirpdZl5QBuuPL
0ieimgZBsGMYRJT729h3usJBgCXz2SB/LC7sMi4QV9yTxcDQ63HKnA5htoPo6yHS9ZBskgldwU1v
B6MADgkKmPvEkEpybE9M7SRqLR+67gUmpG+we7nZO25RWjY7EEYt1xn/pUH/9MYoXA1AdDrgPLlg
Sf5dmx6jv39BVmbvf5jWPE8pkHGMnwY9w6VbvpAl08ZFgHos2NSwr4Khli+dWPaldK0LIx68ZUgp
oLO6vIspYuO7imdZUmvengzaYR0BqkCMTfbDTiz42SWYuxlYMGYVTNVzPopFNJM0h3PgbwwC5LuI
XXoRAGlCAFDGg/6BmGf4SYR8e7aNW3r/Bs1kzjbpGyUw0F9akIkk7AyEAKhxiSFpY6iG0HoLnoxQ
27fwGS0CB4lSkrk3WCpdmihMrseYg4Bru4FngtJAk4zk1MiJGtXD+TovDxOcRb551QvQKg9C5n0T
KVNEr0GeTnqky9+acaAS1x+516etNtlngZiMy2b0e4rn0+k29+joecK04WIeCthXJPXKb1M8zAoF
IK1hXqeMw0q5AD/o68+3FOF7E2a7e4unRePj8nIuDUkhHFmBWFz/0WrJSWWuA8JIbONm4qGsm6ab
lBhHYRtsHu6o7tIxLNqs1Rs0bXRCvSK/+YXevR1wDUcJOLJo/8N0/cN1JmyeZZyKLCe+xh1dmfdm
Zw6Y2XNE0o1dmrbS2kKjC6q5ZBY8cKT25hPey5tTbreqBy0K3YoqFeZ0XvzRXhNEWdIhk9/kBbEo
SQiQybDOoLfovBWVEkHho8pMGCKfEMHo6y6tqxgQq398x3lwH/qreAHF0syYDXkfAaEereiRGb3r
pt3+4QQjO9fJCvJdWIpCAqx8og8iVnoq2fOlIoyZC/IFyea4+J/7bN3ZxgHoS8Z6rYOG7pA+RqEI
2UHTFY6WeeIbcDtoMU1FG4OG3gJBuQwkRLXk/JKfQiUUqN8XOW7EKf/+4B++mtycQU2ylNAxvK5W
tt6hmmzh07YPnNMEyLn0ZVke1uPeI94KWCcs1pMWuVPi4jNtKiDDIUz5E/CrZIAZ26jJUJphVhN/
OCDB3t49W9jvQignULbvD3c+NpjA/9BbjdjvMWwp9LuoKfy2yEk1Kqc2BK/wKlc6M08Nj12GESHU
mIqR6ON8D2hO69mwgjD+zKAjKq055vNAznVtdYYDpYHRpEG2a1T6cT5VgV/2Bk1c17etZzB+Uyt2
S6vIfwnzKJTaW0ThW1LY+8DzqOjHNjnubKVpBmZf6VTMzsIlZKe+qFUvZtBtLX1z9/VX7wQ/BzxK
oeRWBMAczqCf55gQRLDTBr0FTeNCP9AQ9CL3wPwY6Hpmq5TZamcf+2bRkY36TXBjj6L9WFvx3qSB
D9aq9l69f8n4cHCOyDyC+SMOKZYrIDk2Ghqoa7h9c3mznUrHJ2nrHClPAAqOgMP3XGIw87DtbK7C
fsA7hYAp9DqkIt87OxWFQE6D7Ei3azgCw41QrWd87jzW9wZXqVhZAeAuSm3rTUraugXQiB1TIzPx
vfbryp9XrZLSDU6XEV5OhZTbRcIqL0gO4sbdZY9zr/XnifRKIjFuvrpU4dQod5f2Y1pt8EHU5Jjz
3ivBMxASuUUN2MrXW0jxLBvBXE1k3aT5fMxAviviIq5qVoFBG6Dnc4cXiduBX49Lg8ZvzclIlKnd
nllLQUXfcjbW+TG+DjtWOaW+/6J5DZQTyElRriLP9tqfdQi/bjQfvUUajj1mP94pHO76H43Shar7
hcIgMdglR8+j0EAhN7maGhYH6Wr6vmALy8aQtbIXQxX94zj4DwIc+1IrPHStD8VCCdBfuCUH908R
rK58yqSB+jcPf9OFkgKLmfuIB/rOSF7nj8yve4BynPWVF0hHxIM1Jb5dH1OxmEaLvtS2HJE0X/6k
qQlJRW5HJTxqtGSb6goyjRxV1ettKTXkELJRjHI2jDAX61K9pxwGllyLfqfDr1IvNSeGLH5+Q8dc
x0db+DKzWz/JASKMFCN/iQuMs7mFQrXIhT7QmDMJzrxbOe+kCjfsNO1xchTqpLVLk1W6w9N0EQbL
U/UTKoWpLiULlKE4jHLy0daQR4vtsVzy0ew4yI7mhonHfGtIT06OwDEdqwhiCIhJ2BXGYjzLzEPY
D2U52l9Rly7y3lfTeBg7eClynfIvT4MDYKZ145gHTx+7DVxU1pB8D0Ry5lE5pvwLt43P5urmCw/S
MhNr1iWGbL7Ejgcfo4eiBZSZEaD+KhKv+QgYlu+DRiYOD8ehbonD7N63DLrGMhKrILzeYpTMCog7
tXRtn0qWNck67o5nF7uMSQwba3tOE24YxhJli494H3a7Ul4zxHjJLeuRbT+6UU5PB0dXDOQfMiul
SM5bkTRru2PpW7pcXEq8SkuFi8duT3GD4UdUZUnce3pewa/nJ2PmSj7e4O/Dd8CvmwdF3X9XSmOh
jJSdWZ2m78/3dEi6NI8OxsItR3B73Aty//uzmI4YOckp3LcwDV2d48/+XxNlSH4q+bGYUV3r2v40
C92ms2qQjN8KwBPMOHZQ7PIkxZWrDEQOm1TAriCSqTPD2oZktenFKmpqKKYi/gfbbspgViGn3mO8
8YMDg0t7+GX1jLt1SunS7flgZxr2tQsgp8N6zoOBmEDcQ2t3O5AbEPH5qToaf0c5Jc1aQhgA3NsX
zMS23TuwSuk3FWiFuijwRRZUiZaHQD44q/oT8vkPS0CbFMWE0v6tkDnwyfDTGHVXnOAo0FJA7jLn
qpH3tyJIdyutYqyvv2t4Syr8OC92Z6wHoNF3ljq5uVFWjPyI1oSAwbyGLSKKxEdNWaDzHdT/VGuf
PeAb8yDNx6XTd0XdXQbBZh9Kc2HrnoX4LWaSSLGIlBN+udWflswQJXJR81UpS9K1xz+B05YQM8Sm
molAY66Jk3mX7noQsmjix5bv3lD8fZXX7kQMp0Zj0lF8vTkE7hN9h5gPT98mI2tTjsMH78wIQgPk
E48RSQhdyYs9r8qyCvIMqe1nOKpKLM71CXcn/fIxMBm7+LGAizB/TZhPZioLmYoJEPp3FW+2k2Ww
1SxaBw3l9GpzKOfs+Z5bjn5Dw3uFNasFpp6rUXZpC3m0EFTtFKSr/KmRDSd8Mi6AajaVumO6RY+q
SlX23ZmgVaYIq4JsUn1VlplGrK8Cit0DaeeiE5VI49RcoN+55/n0ke3S2I4UV/k9NcCBOBd9IWNL
vj4QW9XH4VH8V/1a0wN3GqvMUdNs7/k4NdOFYt0S7jQ/yj54iWRrlysGT+lK4qL7e9tDARmZD1Qa
ueT68rXBwl0AvvVAKbKEdVQSU7bhM9HKkCyIHO8SURwojBamU0TfbUEiVgWg8ej+Vgw+SuVnUmzh
F1NjLlMTeTZt5YJOQfSbzI+aVzDMeJwcuAM+qOVKQ9CXEEPeA7t0gHQ0KC7YheSywnecnqBsQF/H
SUIjfP4BZ4c7FVietViY/1VfDIwWHVxnBNLLCehC1+lxchUsrHkjryVVvKKkT0JrF9vu4leSuk4h
RmSjdYfiBjl7rjwz+kbhgmEyKDEtgKzhvcReuDloHSQmP9k8GEIsscLUSb5SMOqD+/csrTi0lY87
ihmHPsSwh0Mw/XnWtwzN4mp7gNmMKdKdWO9SDmBD5Yf2ZK9XHU2aERfbUdglXGhMPJJypYjSU8X+
2z2ywXRP4uDbw0GuRztBsjcjzH6jMQ/KTR9OycIBY7dxOLcpj0PM0GMN8RKvRW+Hd1CwBONEQZsP
Q9sWx77JqxdnfYk+oEzB5+mkgDRTbPUMie9l8JulfqI4laJMYCW5cu3b+OBAZSrX8AxUXIkmd3pl
0WKNtNUtmr9AhSO0O9aiHBRvXjqGwWdphSMdiKszfXmTk10U0U8ZiFdWgQKnNPuTNo3aHx64xP1+
ihjeo3WYzisobq5A8bMRTUFTW4RFn0MCfoGR5xJeoCN3TBRX1HKCt9/Fm8uFye2Vw1Y4Ukh+TcW2
rWhrYIJGAeCliDK+u6Vwlv2aWOvjNx4lYWVDgU0nUjJWF2pKXvI7Q0p34nU5FJqsqYvRFtqlnc9c
o265/qNw7vDqiiPdpqZTOv8d1F5dlvWc/p9B83sANLOsO/kvSXuD7KCxev+j9kYVc4P2gs+9mzzY
5tc0IHZ2uentzmxmRTjMef9N+SmCTOR43BhKU89dzIp4v+oCDcqNpxK1P33k3gkLl2SvYT4FH+DH
oS7Y5gtaQ3+F5iYelETYsDn68jKbZBkslz10pAalArcQkMxguyuTDRW0Npowvy6Q5z31I4/2+6nV
DSc3yhbvzRpvP+4NDj0YVc8UaM5CuhG+Tit1hD9DgwPL5VJ89Kjs2LUNy6aOGf53ERvGvU50kW69
5+X6D4gbal6WVz3a27oNEuZsuvaHITKC1UrJ/olGFn63OU2hl5jxZWpWaHYWpXnRr22hw96bZ+3R
yNfmk91inPhbNV68viGJNrRAvCSgnX1vgTtUAzy/sfJefaeVzXJC6jElDD7jsUFo3GuR1ABctzrV
Jr682oNasKeEE74yq9osKQQJ7gabGzmsl7tMjiZi/lRKerpuiD+fiWy5aRZRk5vebWB0+jpHRTXd
Fbof3PNvABKrC0uxCqn6Ftn8GID3NtFqjWUKQm81H301uiYR5N85nR1Qxx48Iduoq8hrdgUchzMF
13MM6PNFiIKgGUXLP2mIJXKyKqcWjEiLSsFlTJej1JW7aQIKNKsTXJNBDXH4PrWJnHxsiZhY+Ikc
8QWJnWhkGmxZ7HwCq2SS9c1tbndnPeBFeUDx2AbKiaqRymNo1KMCScW8SIuAbA6C6h00fmfO5inI
ZXy0KaehvUMwy008YY8+ST+GqboDpeRE3c6PoLbJqGE57sz9tRaIuAShz8QLnYYBi8LKy7fOwlUO
qnmop/E3il+lsWV1ARURYk1P3k6pC0XHKdLxBHQGjiVoGGKK2b7yrmFwpcukRjLFcCV+UTr47lrR
W5wLRSykDqAIQO3xvvOfkx/wDXlc3H4ffJlY66FJn//SzQGS8hqYVgepivIpf0Z+KIzh7pJrLby/
uqgb4Kj7MiGAdq4tAzItriymFYdl2gUbYww8SJqt8De6J8+9XDkTqB0NoRfrD0BEgSgsoRhpitmD
OCFOPzv6LvvXn40XrBdBpd9hvxUkxVsmEe96vYH0mENZLKF71o23/oyltbwhZOIMl+TLoJm8f/0t
mkNYcrhpKxc3zfkg4vfs7qE9fYe3FLvcW1x8/4xO8WcEVVILugH/WLWrLGkbXl0PEP0o32o/q/rs
t8yLiJYv8eXNpBnZXSJ+gapEEz5yJdMrYPyvFp72qkuOmwor97zFDAqhcp55k1roQNyGIqiTQEjk
OAvXTne1X0pOBHzuXDENF3WVvdDsBFFY7iEJKyES0y5HW735qko8WO4NgnzXpLwjaI5Oxavj8TAQ
BNyYy0x2Ppalf390TPJLyANOdhYYUBXHlTemURccE3hl+FHIsJml4l83WMIj9rsocoyiJNHZFdFH
R/LmBzkpiZxvCz2cyviVvVJdXqyN3/X0CkDS7uvZYqu6DGA/SskYwW1I19MZ1TMEc1GYY+McNVXd
2bpsHREsXMOUW/C/t0a3zNjDmr0UFQL/MmOA0Ok/d+zTj9AAlg30cE7jKo+jev4gtU/K/JqIg1Jc
24mrKpHkJSmiDmZjw5FS7NrAh0vdpfi37A9b2AsCBGsaXpBg16okAN5BPwBQu6bK6f98VmPbLDzw
11x+SLASgb3hqcP+eZGYIEVlySm6i5V26Ier2fxj8vEY9R3WdkMN0kqGp520AjYfcWPqES7pCdxM
wa2p5c0Rh/GttsGZPAaGL3l2EM43qeawbqURSgAEBubX4igc/GF7RXaMN7m1O7Ogt+6GSCElxQmf
AGDrkTzz3tu5dyheBX3N9iXc1Srvuz81Szfab9WgeuCPxdImJlaHdVDDKcQfA10xAWxBOmW2kK+M
fLMySCOQbU5hfSauu47ypRRnD4kdrHgGR9uWqS8V55yioUFxA6y9FiCp48A1BD3Q/irAeomV5u9G
6kEz0F/HtshntADEcTjPsWluxCEOzPGYOU5Y71nBAu87+6Oezd+DfCwBt2LrGZzsx1tR/jYgexN9
Hm5twSk+0dzeipr/HnI64yqjWSo9t+QOEugEWj/4crW+P2OB1TZblTejMJYf2Qe6PyAaqfHxD7Uh
MgikgQ4AuqEps59hrhlfjz9vDea8jhq3l3nZwRQEKTk6K6BggPzo1aFMI5f6DPYLXiGn0SMBSD5T
Y8hwfz3kIMcb11fZ86bL1hgJqIzYbAM4rv5ugEgf2CH/CIyGWRohgvx+bI1cnkPwGnaH4urIHqA6
WRe2XiwI7OUaOAMayoKy5Bh9A0vOk3Yo+p1IMJyo0g8M+yyNsMIe6HvfGQFv3j+EcNrkc109ekxo
fyzjr/dGAi5WSCH7KyJpGW4mUutWX0U5NKngPPUmmSs5F5B0trOMuaowwgbk1D1DJouMLqN1UV1j
1OOgWqb6kqO6nPOEjKuP2DUNqkgw4DIK7kHpe2B9/iSiM1tw3Y1eBxmoqZMT7abkTHzumgUXmyqK
XEs84DtnczMisX0IXMD3/nT85yFqdFhhowdbcfkMVnx9PPbp9IFzR1aG8tRZCDP/Tc7mDqGRGj9y
LPsNJrKhLjNBBauKVlaWtfw4Ey9XufzAUAaa62X1xPkN25ZAWs6ePu2fMBcmZleWbzdwlO3k50nD
M3XJ1Bbcx8+eiqg/n3iUD+KP611XnKeUC97YKbDdNJ3Y3R2DVl8DqpihGX+hXdMXsmSC91cUl06e
Pe/qJXBwK5m9+mcI1JwCcN/RTQb4taVag8CoZrXvX0B+9mpEKKJsrV1VPTaaFe2jQdD777BviI/o
rXRhIwDIpzUst+St/eFty7OQwPG/K+WKg8jwjKWLTlUAqvnEgY13YMYqMldSdCMKw4Pi9/A0rpyF
Z+BYN4lvlDTYtwwQlSld+8bIJ8N61RZ4daZKoZ/NYB9ZVEqiNKp3aUdCm9rNBNKkZNT9/rHtdsCo
C3MN4wkeFjXIxmw8MVVBo+3K54h2G/QPLPpVLsXWHk4JSJNR+9N4RW7VQfbGi2EW3R1BOpwcZ7Jv
oKHiJbLp+ytOSmtmWAhCtyeJ+xHkkzfRM0ue84KKdo9i2m35oLPC8Fa93EJ2UN03mHLpVHDrdKa3
rieI9/zq9VQ/tCWG6fwYdIpanqjWkQT6CnrCKa1Udsw2EBXNf1Mm5JNLxx2a0IcpOD/HyZWc4PT5
amP6v8LhOC0F3TzbcmvfuAbdxvt9P4BcTmLWylL3BGbKeOWmxzI+lkdyQEVdnGCdbmzK8jUiXyZo
4ywL2YsbhzdoEEAe/gBWNOxygvc0mpK4g/XaRP2fyc3Z5Ncl+GuKZ3LEX0FHnlFIvG5yRXiq3wd5
k+eMQJvfCIW3Cxrz6FvyrM+BdTlyOY+DzVIUQ+pvoHtjDZHzeppclinZzPPuaWAXLFPQaNiMeGrL
B9D87ngvloAOOPXsIdIzmjYIx5NuzGqDtMXbzxcVrFLuwEBp50DFztXZTC3nTaWsc8khzc7AOTB5
U5cRwIx7dOsIJuBuGvsl4jPYt5iuYZEODkfaHj3mqSQpqXkBO7FdbccP1yTUat/0LZJfwGVGIeAL
CyBsdMF6Xp9WfGHagyrjnRuX1NqtF7tGukUOipMe7zRUzf7pvikdLcWhVsL3KUyiCF3Mn7k95n/l
Oyd2a6r/spieIJi+OrZ3ZJe6fbgzCqcRyg9SCZIqMqMPRTM56UXY+bw+uHUSFY9QnfMAMdyi2+MQ
OeN/CmA2/VSzkLnfTixkC1xUjUdweN5mOpb707BAvvMqUFqz2O38cxEc2r8mu7bthdOL4E8kKccO
oMyO3fVj7DxEIlPHsOx6dUiI5w46VC4au7wPbYgHwlN8u7tCKfTtCFgD4ogSMJbleJLJzUNE4b08
nBG1a1hY76dUgTwW1lj+6KEQoDPRg4IE9CMOErmLGWw7xV5UXyZq/xGqS+rAenf5nFWNu64ClFa/
kDDzP7bRSjM2iZE+bM8eLeAkZ9ecS8KCuRwMaJMy8RQzznt3w9Lkk/ElHiUy0dCfjZ1J2d1WPMOL
I2pbmulrsCIqgp5E8VOARJEvTYGMjg76dd1KDl/cCuK8Vc2/zPoUnA+ZF5+vsyEaimqyvYDD9EPI
6hu+y4Fqh9YyS2bVvtnmXMn9sjqY9Z9IJhx0uakJ2nSHJpK77YKBozXPQIHQ2SHf/XDxV5QrvKZO
PjygO8rScr9rMNqidxeZC1UpfjGq/aCrgrolvg2oGWDpLRAbnZFEJbO1d4SHrkMTusJdTaWfUr3K
tCDWvYdEZmN+t8YIyHh+niHrf6Q9BYDhQImBDDeToH5CxqtPWsos/2cWPmdfTqd8VFya+Euci1cO
rTAKGNDKGkh/OZi7JPFbMB2Nk0zqodOxkIQ4yuEt+Nmz+11PtcfL3ST3GqDA4gI7zdUtf+u+QwN9
sTtHQ7GFqElH278+h68aLPGDrB6ll/L7uvmorA6Is8ncJuKsHmsc1oe0k7bM74r6cNq7+YROasA6
fJX55C8IbK9AkIwSlPbAhic1Oo8gk6pX4M9/raHZV1paRjqyTSw1H6EvrpO4kfELN6CBnofCSKs7
6HbWrutqgJ38+XYB1XEMqF8pf2jImwONq3liwV5rl2IXlp6T1gqnfwODReffQQ2CPtC4lmrrteQP
KSTi7DPDTRT+Qgw4poiumND00GlXbNszekYg2P+ZDmnqnTdIsIOpFDIe/KOObanTxz0fcbi7Nj97
WQfgTuhVAOg4QbbR+X/2IVFSeiEEJkEw8VOckHDJ1Q+hqbioudHcV9b4dEiDFUXRDVT6ENQQjRZP
FHwk2p8BQBiqpFwhdpEhy4MT7FRUVNWhxKJw/ovk6s+iFdlFOTs1rD7IYyRrIZdrMuj+AbAHT624
BtfqbJ6TRYTwwK/cmdmAtT/NaJYwcS3v1aQVphrXycTbVPsav/rwlPIY++tE4WL1wtJ2mtJ4t2U6
ed33lenD1+jU3RyJ3TsnM2TAmltCihMowt+aY8nkt+eqmkkZPlYsvC6Br82zPl9EiBWPe9NB4jEf
vjyz7PG1q8sfJyZ5/T3jR4OvF8MO5Wrl9QXVWGDcqXezMKajVXVIUa6pBSXPFnD2y+3OUlS5vzP8
bQieqk8LbVWTl1Fy6pKo8xHz4ttmjKqbZvDJ6mS8DHsb4JyMTxQCdT4lKsmsqKNjBSCH02a1b3al
lJmvT/yPGz07njiI/uXujMjVixJ73u43DtiRdu4YoqNoD3sq7y6ER3XfF1U8DRUqgDJIFkHro4dg
TtSiMM/Oi6JUuezdnp+JRWKv2zSq+5iI9TVwJSuClmHHZfGpMT1LIDSus3TvhOXM3gOYZjIGgcVz
wcWyhZzZM6hPZBgFHSEoRclrtGXDKnA6dFFcJFP7HTawMSQkcbqtPj+zf8JItUsm1GMsSjqXF71H
3mzQipYhAXdox9WCijl70ctxhX1k7AvkHfkNdMDC4pmR9m+HLS4Iv28rd6CvJIcAVmAHaQuojCrb
Rs3Sx0oe6VicDZ0QNVPRpWSyzLVYngSMKS/oGINYPb6GJWZZJUcMDVwTBiDFboTWUV7JmcGyP3e/
J9OCtHODilucbl4gQMaKyeQ1xl3jT1OvJaA9m2qeycxCc9lT9CnCwsVMFnGWwjmMsgCBQH7CZ9uR
kC6NRyfSuTqpKoOgfskNVpcT1+6e9ErGDrMKoSJpYWUZfXeYLpV8fFBCAxWXF6rQlsD10w9TLrLH
Tjxa/QtYpIKm69r5l33hclCUnk0gErot0GA0FfOwIyQocNSS+GVCFGZZIa+09/paNkrcVRQsmwXA
c3iPL+MqvqfIDDo7Qd+OjofoL5fcfHmr1P08TLT5ILyD8VE0t/8HfbwXJ3K39KXoyPj/aocExnRd
XmonnxckNDHnjdq6MoAB8vgejL4avtWxR+3TudFZWhKpS432ELEVq9Jy4JCIxZ6K/9DrhOfQ1joT
zH+S6HWc346on/i0Eh2mWPbD4Ft/2U3DfamR8c9RWYR+tkSHW9bND8hdLxB3VC+6TCNt+ulaQa29
TfA3sIJaoogtAu39mPkU34OPZSCTiPmv3YfQhnKMoM7TgKJkeopKNkbvqbqjtbxpPnOQxU69cdeA
yAThRF65jyaNQMVmEMpLGByxn5sNHIyP9ENEyi4a05uGSVaPJ/fMQLG7CuJpcePHE0rc2NaDNg8a
5Xe9mI8EIUds/Xnk8VG1sqzLclkKHa3ak/66cDjfGUvJqF0JlyTixZy0t0oOpJLMVajmdg00lMKm
qviLWb/0ooDCJ7hcdhTyG8REos+XSVWenG/0X4MNQLXaHBLd0JW+fGHcWdMJMHWjMX8rGE3n0xpw
FdfpFY0oIKoIKsSHXTzpAkryWyt61k7LTBNjbB/TFaaJttB+fevCZPDie89kEw45MiqIj+esxmK3
ZAC/ffDVm8VC5nz5JOKxZQfwskkLvyogtJlRLqQ4GXqSvJ+oq2NGjLWdoCBjYnjDYk3xrCUjD06K
ldwTLrb6Hs9N+hORxM9IoGyiGoNPvM1f3XL59z/Uy0+odDEKpJkjdLlqaJH5TNpxfiLFXgmm2/GX
9Dvo2DH66tUIwrZntwk7GDJSP1EUtq7JSVUdKxC/Cqbit9i+M+NJt9tgqcJ48LhzqfPyVpQSxs/p
KZc/LR7U9/7lkbX2RMvtJPdhFanF9IeW/h1qnmR86sn50/dzmyqGjlbfceBpSGK1QR5oeffFmidj
J/d5pEa3cn8C8Cy1dQf+sPgfulNl2k2IcF0+BXgksuyBh7EYRrvUvEo+Bv5+DKTcd9H+uFXaVD/S
3Q/eP2DFJgDrhneHog84OARMpF+gTa2eqWH6+9lbb8lW5YmOJxIOS3gB+Jc3AES9NZjHYQEHoiTC
60e9vSpILujU9G2kAXlENRVY0ERGONd/nt8M5meZ7csWyfo/O6mD8ruuZ7Y7VQzkPvP5yely6eGk
AgahyQSOZmpYKJS70XORs/bgJf7q3dgdwObHMRBYmLmJRlVnItJQHgMECcM0/BFWyNSdLpPesHm6
txs3rA688AgAyG1NgG1llmBI/d7JPQ/ACB+2WdvIx3437H3eXfVr3gty92y3VvqVaPZNTY3dJvNZ
LsEb9xGRTh6W6b7l84rkuCBHAHCDmrSemzRhv2UcVOGF7CRqFmlq5nmFnCLNceKXU0SgMiEtXYr9
mtcLqzuJXMHB23u1B0tp8WtItNsvUavONprquwm1UQxSpDn7nwR151odGFrs9SVTWQm76IisubeA
2RAOzSRLftO7AZDChIK0P3icDepzjLjmmOaybIiAehRgOKaDMUKm3vpfsD7KJ6gnqGgGb3m0OTm4
nx9/lk6cbHL+dHeXUys4ocg3BaLq4le2SBE0OZeEHQ5dhY9yUd5sO0nsm/t005ifyKJFr6rXrz0f
uAdQTBCL+COaq65X4FuK853/7EYxxeFEjkDRA82MPGl5gbxlvTHLpUlRMzKC4Z5E6iVP+F/a+TRL
kzHd9JZ99Pz7cyBA9kVu2PNttRlqJFJGJKw2nljpczgRhellpEQcIzHhT0iJO7FDwhilCiDF3Gtz
Q/vHpQot0H/4eMcUpUltzJUwX5oeZrhLh9RtwDohdv/jBAaIrWhSsOWmX5A9CI2YYgyDhSc2oz/a
S40QvZqn+J4Eb+ZLD/Qw/XwdFAPQ+1ZJZIe7FowENe3TVUpWndgr/aE1qJhWGFH8PhcPEe5D6ffx
eH3+55wPx2nbi7UkQgFdjS9golXA6P9CGRkpnedsoYJGg1me3yE8iklJb9K3TRZd2C60s/cOX66c
Ms1SGEGV9q0EuzoAZl0tv6n7RwjMEE9WXZs6M+ztJj3UUH9qD/7lsxkk/RYcZnOkvISMQILpmC+J
9MlMvMIiYYwGoMmd+ch3zzZJeYBlH3AvCdGiWOcBZP+7ZeAyhOq/Y9wA6zWlhISJ9lwW8XI7bvDE
/ts4XZsthNYGtsYtCgyqOl+W8S9D79bcUX6BEDjKYKJdcKgSJxQRZa1VDHZsaVENdeZ1od73n7t8
llkoRHh22pdrpN2nTDrRIGzFsIE+AHUsFKQmRLO9kz1JQIK9CxoTZBo4n15TGOXnW7DhH5EsGxvY
O7sBBO0GlMLi14zOgrvaXUVLLbt1QW5J1PQmGDrq4Oh5rCZ2mTd5FvJvihvDLcRC1WbLACPyIm+P
Ayqy8dHLCpNx5Fal0JglhzPL7l+iqXCegeHNGYnCZkd5exVSNNQSReEyUZmWTdTlwLcStW+gbZzf
C9370ke6bMnGEZ32Sab8I3ti81v1HhxjxeeBwTnW5hyIB4A0Qr42mHiNN6tYVmjVs+9SrVUX6uqE
jgwuk5Z/geAMedWHPE/svAIziF6Yg4EWhgLoYQZdVYHoFENQkNaNX1lCRfL+ABzZGnRV29yEbShA
Sr0FC1E/1c0FI0vRHbgDbPEp61kVMuW83IXX+UCG2m6zw71jpJgIbCNoi3J8wOhvxjHzcrI+Hs+C
LyQJmubyUumAZ76y1ugJYVplwC0S4lDcFGHPKPnk9hsy3kmwhfXkHJWtnHuiNGBi3DBZkSiE9U8k
kF7hZ7NcMzuB7KqsF4eemhE2BuE0pmQsrq6MhyhOqoWXzhkuoY8/aWJzGJFtgS878S3JFRBcuBTC
yzELRXTkP8pKdVz3fsj7kUJI9Ql7oAgnyvR5pnbdDMDpOo2vi3YzUEa0Ii6wVpi3e/+TeNcWo3ij
IrweFi8fcPVC/thb1QmCHx22YRYqGaoVue1SPBZ1Fdatprdawwzy0wPGbuNVG9U9u1PGzJCjEk6M
r2YwuR6b9FVuvfFTFwHHrAyysV5koKokCCuRLdB0sa4HnguRTTiZcQ+7XNptGw2yuD/c5hHtkZIV
TnIj3ZtNTIFUAFlv+ivO8ilyLgXliAK4rHpmcXHiJjvzg1TKFxCx6RCC7S3qxuooRT9bKhbiDkir
RoT9Q94DcmBW3ZrjIznvO6fas56wyX8yTrcg0pjXK6gY4pvl/yR1ZBkSPhaqj3/Y/hN/H4YUMlRd
fikCfdlnpR05bF7V7CNpMjr9AUv03gYiEx8wLQ+G/SlOA8vGkaQy/P5QM/sy0H1gmXSy8U7KdsXR
FMG6sjUZ220ok8rTx5H36nQMlC/hiqnzOmgxNofhUN4bNexGPr9xFy3sG214ZkMj4k1H0MuDTHU2
iLPNDKvdVxGaVC0NqOgkKUCEPNibZAeWJu7iDsqC2Nn2GvQYxEzGza3wXzGHPRCUlJRUQK2SxH0N
Sbf5vxClZk3xp+Lti6Hen5txO9IGJLPyWfWDEh5WYl/HXVoQwWTCDxVQzzs4x0K3qm8WUGZ4sm/H
hlmQvqMOtjhEslgDGaWFVDLHoTc8HuJHjtqER5SJlCdJ9jRAmaKznVVF37Caekz5QN2DhW06ycmJ
9pCzJoSfxWpp8Ud9mJEnDOIRo7kGkvMwmqYy8fNhYoVI63wguDKcLJKv7rSa7QB30IcsyWXiVkeH
pkG5qYvkNA1kqXKTZA7F7QqBW3KjQUUGvL3MZ5+wFqN6R6AaQGQ3h8akyw2oi0A9JrU3csywGiaZ
7q/FRb1OAlypN1SADV1X0Gq7C19ds67k+rFYJvpI1QAVCNl+DeK0bEKboJTOABPfxvZig3qaHeSQ
YbZbsvDU9FAH2AOjDNVlq1/NCQh6U4U4zAcBHsL/ACY1NApxFQj8fpKF3QsPb6KiPvaWx5OTS4Cj
HmlgziYmqeo0XqIv9HIuHdP08GnhzLnUvLqJA2tc9DIdIAD3mQknOwfjGNizvLCUqq0vlq3KGj34
oap6SELCFe9i2p1xww2kj/vp/lDAYAJtKXCKXHKZMUSzqslfA4Rsg10opsVcs21PP4gSb3u00nzz
2XTkHZmYOyI5R1Dv4AeoUrUIous/Mn8eh7B7T6/iYHCcKZnSVrAC4+rrPLVpUtWJXESVxgH1jFGW
S89GvlxI+wwRTHwA2Q1cPBVSzxpfxcaVE/dbzzjwKxSu7E8SnaYmySbgwdhRsSsENj6MvVfAj8el
+YXAy/CCOlHC3N3idPjQB+cbLiI3nGY+Iwv7syilHNjhdKpijHdxzkepkZxqoUJm1nDmFR5A3pau
5hKN4L/rLeig7R/yPoMsTOBEOKIxKDWlO0pQAZI3RvDPPc4gY70kPJFahcWe7KQLwWbNTW8fG18k
9bRsbjQ9EU0z2tl9+AWPBO2uAvvctYZx0nte83+EzRJNHBKdNnazQQlaskELWNJRqsef7L8cTaXG
sNhVwMc6W+oVhQMP6sU8Sm3OOy7LHhDCuS+x4GOybpLBatTaiMwMhaUHNDGzku/p9W03aSn8LpAh
siiREtxR+NiRHdhBwxOe5TOD/Oj+Lu0yGbHyPflqa6a7O4H+GwWkFa07dix60lxxrnsJc3Y+MCN0
xIvSmJK/jDaZCdyPUIASOS9mMzOHimPBRx18wIdJEWcnQoV1vBwP1BdvYF5JeXn5/OIKjZ/ikXwG
96NSL6ANJg5iMvcxiKGkr1zKRi0/Xhz56UV/0NwptV/vK35haJIiEfykhKJU1l/FsKsFGbt4iven
OcI/ghJ8TvABQQoVutRf2G2kIGCUQbX3YCjXLXazOI1PH6Fiwq/7tGvtq43hbUsZvfVy5lVhT/AM
6nAcbXgESJFtiB1ZYd4hW0RiKOBNp4s1bUYIwuJAC4g3W3Ao9j/fd49XA0OlTTo0rnOYdcrX4ezd
6hbbcQ6jE4rwLFaPSZUoEySA+gakViIbnfniZJDFVZsRZXVIHfd34pJ2oESu1gzBoeJ5NRMMTEJw
G2kT0TPLEAI7/TOHSrp24WJiiNexXhKsmuVT9DtlxiKnCC+18Ptd5Q8LY4i9DbjO/O/YPQG2sC9N
h1q04KVY0LbA3bRbwiaOjiAu2aaoVzDX+KrOYABTSpcG00xJFgpWfpwVkL1sSJso4K4yluz1AHZv
k+Q3b/uPy3pzxAGBBDG4Hdgvutg3lcOaxIEIOKVK3p3PkHnivPbYA1h6GAz7+D2Qtc8IwB6WFJxG
fr5V5GDGIGOM7cL48i6kpQUaeJDVikx0X9crg5590VgtUU1XuSI12PacLTjRmzRAwvV5Tpd/Nulc
pruACCWDq4zg+gAsQEfiu832wH2GK9aULk1gyOJe9j+XOWlovmB5O1+cp3iPNLkJKmm+FYqivjDM
TRAWgapJ8iNRlkZ/+Zkj+vlXC1Xq8QnnZB3Nw517O7g+QIf1ODYL/63S0rEZYFQQ+aqa91egca05
LtxzK476Woj6uxY84WC5rjgTHF75vlh/3fQODp6AkkwTTxsPJmPjqMu3M2n3EauX4qb2YVcF0q1t
11u4rUOweKrqtNrhpRMnjW/GWASIpfpj3BrXTRV2JG4tw1lMCYwV/VWk52Y+euo1fWMi9Dc5dTkC
2Hu5w/askUfUmjsnwp7i9qs/FLG0xw1U5bTSqUlsZr2XHTkO1S2FCfFq7u+uZOFWer9r4VL+CG/C
rFPsvjg9GtM93a8x7ygGcF51Ogq9GoYPqfQvx1tbwWC49119pKTVfMy53JKznaRx8mlIbjH6cUUD
1uQyxc4WazOeOA0Ds+LqaG9oFFE/QGwrSyPbSCROz0VW7LPrrzK1Z2QPr1SoI5i2o9c8ZClPwKMa
TNMAniUIGJkAasPOXa2y8mOwrnurEJ76zHXBI5wn0yh6Ybg5+nX3MKWXDbYntHp/hPlz7u3YfPQp
PNY3AnQqh4bluTyMHcLRMvxFNkaEvrNW/GsiakhqKfalmQnpo3YgrKEcmvcBMbVChsCWQOgjuOcf
s80H6WzJzUFpbOx1qWe89WhTePxyESuy1bDaIL3K/rQtNhoIUocx+zNu+Kf5BsKycgcQbIeXut/P
59X8JTxpMabUCym20R8JIC+G/BZmDy1rIbIJ6ll6E7Fz+6Tib6s4EHpYzbRYe6LlMVjpWdEU0KPv
3AhqBLQWAR2MGUzLXD1ULGxW3fAdmiuA1aVLpUk4t/mrgpL2rs2fn7edipGtnnydeGlbxP4tnPgi
OUmyfkYPKnV9sCOW9rZYHqjJfxeOI6Pk0PHGwZaMCfDRK8h96Q5qNXKfDYinMUPG2MVMRGbvOSsG
ikfPjLcmrnhZTEkjiydvAFyAyo5YY9sUuqZ8W4I5qDvUf/2WiR/3GOPLRbB0j9B6ndwJegx/Ggkk
d2Gg09lCxIVWFpbGPQQIxuklQvvFA+HOXj7A75NqC7f0MiLRmmpY5WeTGKxXBlKHExDzlqJYf3vL
Wg2WZt9YYhcqUSFoyiKZ8UslcmFar6gquOW7DXGAjMB7aUasmKjpgXWnJLNIgM1eY9Xav8T/q+on
EqcZp+/pQjbE6d9Pqcul+uy4JSPgIHPLXZaFA+GlHs1lDxokObBUecNgK7lrbgWLBcKywSnk9TVi
AC0glwoXDJkFqlB1LbuwvQYXk2RGuV6N/sOh7sHZX5b7XTdCQx3l6Ki0AXN5ubNLTIIQz5arlSZE
ReaWJZbGFu3lae2Xl5wmqjSJfiN6kvrXpiY0MalzqAqxp4XXbh+0x9qhW4+IH1h6Ok3kDiUjS1Ef
q5L4Lg53q073+h3ZnrGp6QxMuPiavUvxyAevWZxka1Ewxl2s+G0LW7tVWObe1dAtv13ObbEFRB0W
XdEJ5SqWgJTJWb15is9+09iIEZe5J3n3SQrG483YsuvuYTZNqGRjxt+X+SN2kXjQhLfEzF7urumQ
tDnk6ooouniDtvV5XaTGbaxSvCnK5I2RDKL36JJddWVYP5xbMQXneG4VDZZjmuqxUJl/RoBzBXQs
NsNiiOeYFT9xDWYPNQ+iNQ+8/JJOEdaxRgOJwtEppWgCB/7PiXRxmnrS6gtzbBC/oqGV3aCVUPVQ
rfNyD9mTW0ljYxqDZyTyLiyHiu7xt+zmTQHWuiyicgq1Kq9BGKKg0LdOM72SC8sKgO677DeYHLLY
MoOt7HlrZSDDWw2WJh2K5sPLJgQqXKtG2/PFjx2xTrLkP2qWhoLAfTLS0nNXabbdrOG+p9YtbKY7
D3l22f7pkjzBwTPIbqKi0GNo3zdsE73Zsx9W+6G9b18MHKjSUpgy+Jdy9fxouadX+7hC9OxDLQsg
Rl/77za4D6VNhMVctz6qs2rSrRZQpF+nT/Zu96N8g4DBEaijYrHzSgW/Cf5/P98x4SLLZbHQ2rbw
TBsHj3OoxlnNech2Gpa4TDGhbT3fuzRv6BVTQbkb+9kkussEbdK6olOmZaxlq6Ap2JT9hSrTd2Zu
VWi1gFDW7WrdWSNIMzTp7+uNpkIx7yq9p64gmIsej9rrFvj/CFxgW37smcDxHEWtOpCw2mKmYkaN
VMIBaK2DgGYgMEPLmQqdI9DFpY3q1FoGHmHvrvppPPwwmNSA6S2vY9R5l9dyuXGEoVfWcTqMCZOs
YlO3Em0V50pfVxlNhv9Ws7JwDzTVcxYt5ioK3KzgKrSWn0RcrC61zhkTYNEgeOm98dLumtRAEE/y
nl5Vsii/U4Q0NuHsD1i23sywkiUShFDVtsBsRyFXLyz3ebvgSFNJH2+MLlFnyLnsWTqNJGGzBQZZ
P6AJ43PJxmUT+G4uySVei+LAS2rv4FOWZLK2qfEYZQuwnq3KJaZxrFDQasjiPp1b9fKDNlpi7hnq
Oh4himy16vIaPurlVPi44xmAy4GQB4nCy++nObesMY0zY9BDREs0dq88Yf+9Hz/TARvRhQDDeEzX
LZWsUt/Ixl8f5d9yxeg5ERJlALJmfuvAd9gBNIRy5spK5XW/ePpb4mIJF0/8IyVoaJMwGefePXHu
CUmKS6qeTgNfV5iF2IKnPwCO2gg+JDqSBwYpThjFgUR/PiPcQfNgtBh/bRMC2XgcgV/13rYvZLmC
3eNoSMoUGHtpiSRDXVFFORjEJP4ZnKcAz1tNw7C1vwLfAhyRbqobdofKjt184+R2JHhRxyfxSKZt
f03n0vQf2EOlqJa/ThlQTAAi2Mr+K026MS13UuVPMHAwzOUiAo4rbOjwBDKnx7wLNd2nqx4COx++
2UUok1cfIvpJj4rtG3FvdDZ+CeZOwemSZzpuMgzfWqmGLR1/fv+pFfEwOMajOVBYVbQh4hCSddrh
mECaeV0wrcNtuu2hTeKq4EhaKXlntOIssiYCnapbaIYHyHSuKqZHMN9kvlaU48ZLMaUlT3NHIcct
JeXs3E/UkBnm2cesaknmQIzATTNBGSkHQXAdc9bFhfxJJbMrLGv44j/4MitjaEF0ugv2bw/Zmh4i
YAsWmGQ1vgehHNold5g/DNB6kwpjRsRfeoTHOX63I/Bx4/iP+0JOIdrFtGY72Vk8WaOp066+ov5R
uOBWeoOq7eTqS+DFMSqg3TXtXIN3TccqCUVRh3BtH4b4i5LsXRQW4y7FQtHcODpZoqt8SatkkCLY
8y/5d3Xyah1v4aUhpBBgJjzJtf4r+tWLDuNd34TITzp/QpqnvAiUnn1YB+2e+TC8fxGtGBAm2188
r3DSF63/Lr/ILMzeRqYc5DTzTp43Pg81U6ONk7F1K04fvvhJZw56OCp0gYEOaR9rtC3OiYBMedBE
dmFuCrj20k5785jBumKgcSF2M0lBieEbtHo4pzCp5dlh0zgrECWL25Ha22Ld22tsh4I21mhJgGB0
jtUMWXoQDTkEMZoxlKBdMIXe6I6xbgEZE53XPwJAKqGbALoMQIj2l/NJlBWtO1QIjTZbEWXUoUiV
DHCR8fFotTC1XkvH1Mo0ZelvMbIgXe58/0a0zLu8vAFihwrn32r+zt1XqM6MSAV6xUyFTIX25zXo
OMwopWTfyU1rEdITF7LlKhSpAD1KiBMIZscORVgyTdtVoz2bTRkMmbn86iYULVmMAcJjwS3mobAQ
gMciY/CGYMf0jmQvf9/OW0dzvnId6o6XHGQ4AylI9XUVfseO+dHLzoqTM3q1nnqt/KSplDqHi3Yg
xujkIJ34KtaSKhsxkiey1sN3vJbUFdRxbObAaQWICnvnfcBJ5y/QE4NE4kE+EUWqLaxycRBnMPnu
Oe2ppBsjmT/5dLuRAUBDr0YCveH4Os3lISmI2xvzGbCF8+NaC8WzjSazCIXPCzyoXh6qOkuzCIfR
w4KHADN2xi45+dsSG4gnN6HrGRztyl57Rq5W6nIOsTJigm1yWfASiTO3VLcMnpikVPSDAPvSeub8
mh45MsY4SIgZfGibyeSwhqUVxj3/mylBeJYJ5QZTyT/yU/eUwuaIDeM6i1d1XEYMlHG4AykW8W06
TvBt7MJ62VN9ECWNbZRaKhmWC7cJ596vsBQfCiDcRTW5pOkvTLryZ5Tn8NK9RzQk3Hur6xI8pywI
k0q8Q1+TE9eW1sB3oxwYJt/HF4iraXkY9fjs1k6pi6WsKMcPVJXWLCIZIxS+ggCKHcfye/dPsbXT
ZfllA71WSaF03pNdjLw4ClGl7xcXx6CSvBlla9EEwhaOA8b898navxZxzv98jHdlThaA4mupHqw1
Qw0FBDc5K7Dvp3Jvd+wyHRAIQTHk/p004MMI4E9ud8cbAW8gpYY36OZfOnYc/K03tWHqVjupt0hH
BF1aH33Y9ES798Q/9JPTlKjMTXR28apMFlmWaAs8zO+ZkFhOhMDkj55/eHD9Ts1E/RBSeB71HktC
TLQruoFoKsZ6h2kvZFsOvOAWG/VFbsBEmxJjgp4Nt1kWYoW5PlV2nhUAj07NDYAqZpVVykTF8a8X
uuBEBg0c0HtLK5aN3LcFInNfRZYZPEPFNlRhe0YyCC/UIGukKIGJ8ZmGRXw6uCce2MlZC1aHCsj+
CjCouA9i6N6ZRO5Mb4XNVF5pZojC1zMxx6FHeKNzEQNXX/gvIASkK9Ir9Ggy7RvXsp3t4G/3aq/5
sjqzC7nTOWC50Jt/YTm1Aikg54eEnM/R/nRe+2G0wIMbPQOp9Sqh2T50NiNYB7jjckADN7z0K5MV
SOAE2pn8TDztpvdwPnFcb2kTi1qqPoZbMH5plAkQN+01UOQ/zx6rXk4tqxXm5LaAeBTNFXL466eG
SCG2DW49zTCsmCXBBC7UhIBeVhUd5pb1jbtx7ehuhhwbSODzOnyD/awiDYEXzamtWZbn3/IuGsL1
4LFtjRn/FYYjOcawRHRH6IZpfpAlg9kqzT0QkxlNv2E4+9rGDDXhFRrOr2gNVf2TR4ByknwGbVJe
cYAqQGaAUY+duJvjMpZiOS23ZU+XfAJ+Kl4BgUf9L+vlyadJuDO/mKwuDMsDEA243afGSHv0O7KR
x9UOUIqZe68d93g4vtkxF6Ufno9U1SvqWyeTybuF72/2sop6Wjtq4FKOC0gnjVy0dmQtNd6oPOUl
V6Jc6VHe4a9zKMgTmAl7Pdi9pSBKXhjYBOqOUyMOlGh1u7b9ZOZyBy9PQRtkO+uhWqmLyOtwSCE1
Sde/A1IfJZ7jS0VwwiKM9yRjMfHP5QQDK18JFIIO+azOOy5CntCc90ohdq7efYSB/IR3HQGWqq0S
vZsARe6cUAYiH8Xvx+lX1KQT40qixixFt3xamIlqSn6tDkNegxSvklz9VI5vLcytKZIsxNBOrlDj
Llfuh2X6ODuX//YzANzAWkFV0NNmxnWaAOtJNyOaiEc4usYTrUUS98WjzpeZiiHpQ2AaDdoTiHHD
tn9ftVy2hlXY5S2/uZVP/DmltAnNH1RjrpDQAT/Vwki3sy9HpriLxxXZK9P4bXZFUUZmFeEQM8/i
LhZZD/SVmwefmhCUvTBEFfM50OVK/41lzPj7N2M92M51Yx5tK7DhRwrqbrKgyRHpN5rI+bUljJOU
0tVRimwU7iP2SRZQWCfIhGjpfHIvARPVQ3DMftjAOmrnStS1NPlLQTL80L4YehuMB7S0CNpTgEem
Rm/l3cIRijVQ/8q9YZsqcjbNgQfLYz7aJPrK351A7sbifeTSc5DGo5s+Ei9hpPeLg337sW45zKJ9
lqHLBQkehVLOiW23O+yvZon52YJPTQjlRfgSgD+V3CTsAYjsIA+K7bwfd5QBLxG9EkOo0ww/gy/G
qb/SJpxtjx04pIHISEvhEXFj64vEWXh7xrycalJtWBGtsoN9u/I//ClMizz0mM3Uxc5/ezBDag9e
TFASOk3AJzr+JdKh+P6DVPKODqJXmiDz+xnsybA6oDOypv5S9usafunPXv4mKv8K1Lq7teGo+due
BEJGuCL8WQFMMKAe/1SGVxRnoMQW0CGoC4kvfeumSDUWAmig0V/UoaNOSLiriulm12ubgaRclDMa
Y0TA4lxlR+NRK4v1HxnWtlvBLLV1o+20TUlu1cWEYW9Igp+VL5Eri3HSgSOWMC8y9FtpQwecVwhi
riE1k5g1Rw6u9ZZauQAvo6FD7dLh8mnjMLDrdruZaS3lfPGqISaWyWLu+Sv33h1dHbcJZhi1v9wM
N8kPVgzGE9s9NlcqqSUUgu2QNNAfjsHu7+e54KUYofPVsMyBk0qbUMV+/oroaWM74SrTaIcq1wlT
wDL+VzvOutGm9DBnlrZPBGJ29OZ5t1NHtPOezVCpevGfVB8S8cYUuOyu42mVxWJLrNZTN87rns/p
WCsLmucm2idegKxMdea83xZPGtN4v+G/Zkh1EUcZbnu9G3Vja55xpLPdT7SDaim7DNlAcW+eMi6s
X7azvJzNJAaKjDdHWlaNzP/nSXlR6gdg2XrGSlABjmCblOt85HyYW4CRfxCO1BKaWfMiqfKAwb1r
Wso2EFnAEKd/BQbBBS694rXPZYEiA1jiHveNn+njqTZrC8IlBFi1DkojHeScYIF9XFgqm977itGH
mKqdF5uVSZyiORdeomiqL3AYagH8TDnWDMWrljVRck5zXzn+yaocVYgEsxKRXjMRbDnRr2TtfDkQ
E3KGqLUnR+KxMDtW15Sm4VCYzt/0WnW+oX5PRQ9x7+iQ83uD2JIvRXs4BHlU+CtPWF2dKb9KBiDz
zg2jC5s1UWPhyYLyeVDZkzWRugmZENHCeupQDDk4vP0KKEQ1yRj9XcqEfUVbhP1sDbMpta+LMJ/j
4JD0VGqkkE7L/yXbCkukrWw3YH0xX85LP6M+bbkzzAPxTQZ+KMpjp/vuxUP5wZFKFdtIDCQfpdLi
R3A1KWVJBaDVErwSWhGx0fSx4wng0STN6v/TAy9X2FYGDnvkx76Ts5blMGLOm/0Yl5S+Z4paHqdG
M5eOmgEJ5YS+Til8qPlp5XKk9Bs2bSgsqe/ARTbt4lz4y6j5yLEJD1k6Lx/RfLSydg/rpvLgV2a+
/Wm+f8EQ890X4tB2WtWBfq8bscfbc59L8djjyfhxv8vxzJckqjUMUouAQB6ciL/HcWR0bPcy58Iq
yE9afeum7MdUQb7VB82DK4nj9QK/wsSaxTf4AEtsfXesdcvp6AFfNGAzxIaLuM0os3uIlLRaNzXo
zxVjUOusKXNTmpdd+rNDH+OqwXwV/E4ZRVy4Ukjtt1m6tgCePZUKvlgWpGxmP1X8jU8T7/F9lPb4
wb481+25NS7UY8evZdfhO2DjZARzUrxRK2Go3TW2v90ezRBoaFJuh15YnwBM1QlzzVQyly3N3kBZ
48N7gzYMfoGFCs0GgfnnXexbGfibe5F3gUka3Eqv99/EfonYil48c1+1LwsAnbhOndo1lOd4cHJ0
6ibo1P/12LjLMoGDhCNzfBkusRvFnaVb/gENpk2GnTFe3lx1E8K877OCyi8gThgiL8cL2tWju/o1
YPLhp8rf/Vii8NWj91nltvCgynDD1aPJhNg2du3f4TPZ+vzgWUzcbH+52E6lhAo9SpzTYU8e+o/7
NJobznvCvmNBe/iObk+klGjgazVomAWfaiVO4Mvqlde67uDyZ+bnz8Tdt5zYvstSjc3YKx4k4FF3
boJ9341oOgfvZJFNyAbS0HvFyDB9E6WWayZE4lxg/Gwx7+IqOF6zPW6lUVmXtDdmoSjPQy3QBqly
MmiRg/yAs8ztjJvHlrHVtafHwN2kiibkS6v+snD9Bxkb4BUi1yDWa6xp9Idouvl6C+rFzCR/6zY3
tLodAP++WF1kXunUdo13SZbRvruWw6AmZCB+sY3KBQtvVfUFC2kokrCfk1AWGrQ1YZ+JPUGdnHw6
n+Dti7lk4uDdkoe37pLU2c+23MBjPXikLUwPyXOX9g/ms9mUnTm4KmCVmFOtq0nKedExjcz2DbgZ
7XXLcbPxT5Ycjyxbw1o5f9lL/eAofOJCrJAJbMYVR8aj1Fn1v/2gK4zwt9oGK9IW11KCR8ZQWk2W
k3EieuUC6jaXG5U0jhXRMmHnrG++VoIGtxnqjD2dkb5kHY65A7f7P9z6oWX03SKX1UPLn8jNc5SL
pT3bjZRg8yRgnpHds28bdWxQgHrPFhWwL0hMv4FFLPvii0rjEJcEGuBAlCEKE3XXGXeNbOmGrxlD
DxuRsPSerIVZxB8Hhspms5xl/ersFzq8hnFRuXsI35IRzqDlu/ENWcGwHAMNfNhaAfeuiIAetM3k
cTPq2MKmuhfh0JHzHDAGwnNK+PTpia5i/PEkd3MiW+h6SUmF/AxDEf7kl4RvXW0VL+XS7oszVzJY
9K5GZ5Vhg12OWPAYWrZgAK8RTbuYk3/kwTsynzCCXHvVI8Zw8JeIdOi/SvJVpHqTcVJRW9aizR5Z
sf4U5DrCXU0/Rd1ttaE+MHPhnDliN0CN5laA+ylWrKdY8ivZ5gjOHFoup6Y3JrXzyCt3S4pDzNBj
QJKpWA2wkEXedCaD7thbpp/6RmQUdt6jxYziCuVXOrOVq/VVwiPiK5YLg6NOSVekQA4Zw6mVWE6o
DKLAUqslRw9SGVIShBXedpyjvLTaoeZgyx0D1GAOg+1kC8jZOy5WZwUJET1hFDwVbfm8azeJLrXg
142IGFhnMJ16lV3RoVWh2a4v+LwQ+vMXkc3HvVo8ew2JtGKKfeL5sa29aW4hF3bZ7rrnmHcWtzC/
ZkegjZzbvAGuqXyH5nnzlLv+AcT4oB0GdWquN8A8yYdem62C9W+pN0wSKi0UhrXgvjdXyy3DjLZF
A/q+ZACxZBlHoThYoi182X4sRJ/fNgamX2HmrLveNQA9lPESdMBk84qOcXeOG9EGQ26fz/2ODGYt
peGNgbwfkGCWauNr6eZA/t0Qo+UC+ouCEHsY8B0uSEQxEtbRlDsh+huukzSUFe/dz/V9iSlGQEcR
M9Bx4cd3Vb1MZDS0xKqmMItmXAAt+W80t00BRRAIzZ2hyvJ7o6Z5DcuqbRv9ON3WIsaiCEB89PPu
8BDtqiBnTtolrA7mmzK/HAo6Dq+vjQF1l056QfdFeF82fbJE/cLFpKyraY+KIQ1U+Hlkp+dn69wN
4ckMI1M70As4j4XLXG/KubmLG0A1j2/f/Y75bK62nb04gRA5XgiRK4eICgMc3cYGW1SKwNmDCo0w
LoaglVXxfPFKS+Vrk4Ox336s/kAHA64JPhGhp/a+GXEzw+wspWueYL0R8JEi9Nn1kYLCSHfuBZm0
9gMrUfdbJBhBQsTaAU5Xq40C5eHebeOxS+KAUZ/jh1bAKfS/tRupuJBbboQQNAAk0QXLND/XejWM
uoBiAwgiycCU17I+oMd7itV/qfTR1GB1+dDFu8QCOxq0xvVZVTjEMizMPfQfIFZKnrEZ+A+tkE/w
a40IOj/ZTaDgEgLtdAm09EnrDGcROYX8mDPGd//tDY3cynDwHfsmDUwPkB7DARq8cvmtQxtLqwIO
uUN/Mk7s2zUIPstZWj5S35rWGOcDIXJSLOBmM8PAfIG4rPZf3rSoMxqIshA+5I5Jkpfyb65HpLfO
TV/ssgp+PUKz+nrAZYpqSSr/4JCZdfSCEaoYtnZJTjlt7p4uxecX0uoRn6DoTMieN73bfkfI73VB
DDYgRwb8m4mUIqWRaLQrLoTpd5kOUuezbtZLk2SC68OlfFaM3W+UqTcgQ0IcWgnB1jkbn5712PYC
O5yyYONvi1AenDoepl53dmcjHII4ya37O921ln/56GQWGj/j3GAbbcs2t3N/vLEUOULyG5JlAK09
frTWoQEVII/gbMW/NXxgqBn5nbKRw1Glt2KuNgBy2r4s4IZU8v9VheqAoKy3X9YQM/Gc80ODAw28
rAPhND8AgYaZ2fs5rTKSV8LnHg9ju6RqeXvngue4uskI5RzLGgcbXkAE0D+powGZZyagH1eE7KT0
3ORe4QRipzi2RZ2LX0qTTR+/Ljfc/YcD/TATDmtVl8FTveXTqU/bs3v3thoWiHgDmkpPwv1ViQZJ
QN59TtvJ43vyctEyYmhlifrzyQT+NUksbaPnsD7v0T9RvpGoTt8uIOxLnAYREtotg7d+mFIeWCfx
28uDOn30jfBC/UfG1PzQslizvZ/wCipQI56wK9Cs9tHpLwnnc6m1cWiZaJpLleHzPk1ivt+z+F+G
ZUh/mMaPIIKQix2TlN9liUggxzTgbz7AIRozPe3G8rhSdZBZ2F3jaH5Y/GonYkx2RWJ0i5pMl+XE
xINiOzprqyffmHXYkWNmtR+qPVf5bqNAWed71iG2ZwbmwomnvTHCV6qaqrA2YVozyoEqZoMXiEtF
cCwVMyu/t0SeJwGZR3H/RmIfbHD1krRvBtuBwlcyP91h0PGzOorgBqE0V4YNdG9wpG41tvxiuv91
8v+KIN8dpsFDJ/3WE0PonjkdOg/m5rWQJVVar6HRwLmeIw5KxNab6hoiUcrE7U1vBRYuiddAS8TV
vCOApYSH5fnZmvcPd7NCqilo4HtKUzunxDCpG2ArA8tufFWZKM7rlPkYdWTeZA5W4Vkwrua3+Ns2
p7bUiBsVEocWtXe5Nx/FkCt4NGzdwe2x12PhHqaC8Pe/bmWpWt3wSamMQmB7zkfw7yJTvE5hIooH
gZXMCQZh14ewAtnBhZE8j1boGNbLqb4htUfkEMw1QB7KSsDKfgK2sxVSu8ErT9yR1QfiqAzyBjVr
ikt+ky2FyIMEvyKxsUK8C1DWtHSmacLH47WzMbqCrx9CVra30i/Kwms0yqOOpkSC0mvBkYywYSk2
Z4IqMmuiIc743OsImPsJIVeCuCBc4sU7lrLtgsk+pY6jJWjVsN70kYRt6r9E0Drgo2qs5ANqvkEn
ofmqSAkfyIpLL1x6pU4NF/y/rzwEQNR6wR+LuzCWLgluvK2xld110pbhXv2A57byISOz3PlexQ0x
QNcbCkKvZoJlAvqPsqrsp/kckgOZdagjWddcaTO7Yh9vefFn+FmN9S1B+PAX7xqZXMcjZ5On9n4F
cdjDCzTF1hy85ljHf6CoQEx7T0vd8A02h1FzZN+jtr9flmSIOifoqDmIbi8iaP9EMf8/JInU6oVh
YrmWUysWnigIpfOh7EUO8Mbe2oLlRxmZpk4aGca+41RI5dz6aeHeP00295Yzn7AJbRhcL3D9W5fF
UzwalwCWbE7RYvAazwJLlEqfrBc031Xsq+izc0BLqRAJY0c3FH1H9/PDTRViL0svtiPgIRwtp6Lc
SdLnCXn22fUeMd2SuA6LNNUVYU1Ae46IT+W8cMgjpYVbUnfOs4UmPzERV3GqRtB2D9WbhT8I9c5l
+2OEl0yXmufcPcFx9o0GfNo+/uo2xQKxldzFZxJPrbB6uZ+ADTe/lg9e3/T3QOPcJqf687Y83ZX4
grCcZgciw4euO841W+qufOig9uDRY4omrjGrpw7pYsOqYnYt7kD4mN4z2aqGjfzT/rmkmMgXsvKx
kySY3zHVL59u7S6DhmWAETO4wmS8eSoK7jmH3m3t44K4w16pYOGUw8dXSfVhLwOG0lFQcMiK7iPX
1kPu39dRiahwkrOwGfiO8mf8i/RqJy+CQ0+68cXGXygb8lr0O4NXtOF99M+dzcnCdJIGrux3rM/U
J8gKszUXhZf9BscI/TFjqGcvP9Yz8LKRgd4n9Tj47vHpSve/ERx9pQ/92lQgtnc+R9aot9LfQV66
yzjoRlkQTKDUJGNXnL235Tiq0H3fCN9t/7NLoF06QT18CADrGCaqjjrzBWXtBtDLm9kP1Jm9QwI3
XEhvrOewGagX8Rv+5uzdGHBxsk8v5K/KC/7X7zgECq1FolnsW37t0KRGClOqEqD2Y0ckUMZzFe1K
bTF6MWpGBgG0Gr1SdSi8Y+Vp9L4leb14XAaKNXygr3dKkperQFfMRm5KZyXXmacWJtSrEEOXJBL+
7MTOBi6AElIehQCq8vCSgxy3DTsXvc/+dJkNh0BbjeWHqiWUWi7kFCeFmcjpBQa1byVvu5k3o1ub
wAPoarzWcaHjCxWLQDZS7S7wAr3rcaMRiz0uaeZyGwgk2+Y+4fyrjugavRLWwXaqj0+j4TuiMOK8
RCN/zYj7g4GLX2nSzVxjPUmch0k29ai98BWrn9hb60SyEinu4Vdhhyf8FTjg09oRvoNJqheYpPi1
KKKcSXCyhl8Z1Ml3Eqh6kWKhOxCbtQuQtzoPx9AttPIRgxV+HOQmfMmEmQ3feLVbrfV9ZVUBigqU
L/gwNg2tA8a3iaeieCwm4OKNahLJADoAIAUoF+dCsV8OIubur1jIavoCa7GiKOP9KyTGSaGbuVtq
iSUSp5Qv6M276OtcG7tUSb4tFPiYmI826Xh2FlrH2kWWWYh9Kf3vML0z84smAUuEAghQgOYia7t0
M83fBuynC2lQHU9YT41XGFB34YVIXIMq1keePhWeDe+VQo1AGg8uaF3gRMnbqVYIFrXjAPHErfk5
Rz9LsKWO0xbpI6mYGTtxs504NUl7xLweevJqXhmL6HD3oZP5/QwVNrYLoVFP7X0uFMNnnelQFWrC
oX5nIPQQgi3sYiu6Gw1VCLIqWklEYaf6BX5+Q1iV5hNT4kah02eAXsxfCtQsZHA9aBneBhUNhy29
id8WalFBlknyMP2jHI3OSCe3vrlKkKqq9YJY3HVO8gPWpXQN1MmRPRa8MyztXaOWqTD2oBRgq3El
uNaQrhYuS90c4dDcv94NBbeaJ/ufqyVavVcGCA//X7buNjNDARcaaFeKW+pJhlz9U0eNWzF0jOw9
7uTYIfFnW3Wf6mTAQnikOE8yP6sK4mX4mgBfaBd7GeiBGO7CHZHROPd8kiKp0ZIx4Tzvt5LMfceK
y4kUP1A2MeogOe/5ZVdQ7qGxd1X062e6ts0Lsb42ddOE7fhNiMK1Qdg1FvbCOlqLX7LGYBkoVGmO
zXw6zyFSyVjvWQcaxmSLESKjvSJTKOB3nqPk0Q9rzQZ866iJ0BP8gusvc5xI51TOVsJD9D9nXbBE
uk/lrUyd41R6bGCyt6D3dg5x9TnqtVcmdKojREKos7E9j+56tycknblCozdi6hjfD0Xm2VL+iv6N
p8ryGE3RuZ4eSElcY02pZXCBa48tUN+HapCL4JyhRH9LSjAaXJfK6lA0s1uB+wf/DYgsFcHj3TVh
LMAv9BkwDMXfnaUyyPauZiyJ309bdUaQWvUBEzUaOs5M/EC8tRADm2VqHJp2rEV5g2NeptPmWZvw
JyB5Cz2ddK3Dkwh6aPoFzlxelV56Z3tqOIKPc1jKq8fvMW7g2/FivX7/p3aQi45I5aPe24K8vfho
R6TGvRCWGoytW35UXpEjB6iubiRVrH3OaEujgvhyVPCmEQLdL0w8AKix8qaPPgUX7UuuROEGgo9N
9wfsrHp7U7dha99F4QSMP/glnVSyKZUj8MdUoRHPARjzV5GLTayyRwdFjqa4JRro65btJYAyZG0B
b4B+mkHqS4je3/1p2jcX2sRcSGCbFCb5zQ4ZFhhZ4toMN2LhXD2acP3Osm4GKLC/tfd+l/TNHRBz
BLido+zyDnznN9bH2zXSmLG7xSv/ZEmKYYoFIzMBfeDNZZ6iviC47T2S2yRa4uGX8TpjIKjplOa7
2cGmjflRQGQ+rUQ2O7xJrWqloxocuDN1lyUPqQmnk45jHu9ViatB42bzn7KzovqhtWr2rTfHRf66
s6PrWVOPe/HXgJTHlqihn7Hty61oINUB6FVD+TbWKxHI/bZDpicj6gMTx7ezZMt4KYe7zT6IsB20
Em3R6LlNAP2f9gH7iaQPJIqLbjMhU7O8P5p6zCMgZo9gHL7pxmeGkdzdac6eKeEIRboumzeIDiZi
7OLvyak9zto3Z2hxZN1r7835yHBW3XlN2BrrKTs9fcjU1s870XS/yeMyzrn8c2rU+90S+tIaZH9j
MTQkPTKTaUZaWVWoYPTBiB5FRZ/hJRxbq0DyMcySDWvFG+uhxC6K3o1NxUg0FpF6mOY7nOEDVKy5
R6Zonu/9GERJhfAO79oCwWl8vGu8IKKxCDf8TMYLuwC0umBrp3t3KuQOQiLzQ+M1zFJOXz0SO5ZI
2XqVucXgULv1t4ggeMvvhEo9t+f7JYwz+/WHxDv1LFz83ihhiy4ODlYTsLH1zykdIMAk7vjspBl5
VNsB1hsIWkGAfHCWlVYZp324G4zEni52vPvdUbXrAwYg8lCSPg0UvMYGTYKbgh74FqjuyF3tCv2J
FZVjQ7xD5u04PsNj1MYpEKU1bhy+hZZ0GbtYGUU9RF8VmkFxASamtXcT1ShP6tFJWDIz0HSt0UvN
G5lyUkmOEM4qOA2QtUGiCxiOAxXNIWFlL91Od4w0kRYGTzMRThRz9jEFREz5L1ZjIB3y/b/F/uBl
z1yIqFbE6DmUlmbK0W6kNgYYlh0GfAa6i95xwo7GwzzQL86MClU29rpTmLlCDU7iqEZ8NpsBPiSV
k6afgCvyHACXpaX/KfHnxPr8SyCw/LFpfFTR6sQFwrUzXbBDFAKcw5yDVFJfhqLidiknDUziaGN4
sL/NnhgZ8wIbiVL/trH1TbGsJT3xkzrThKd1trklnhHMcwzwhmmx5OOGhfHjez1HyJdwyezvPyKZ
TIfOMbmM5QRnr82Xiw4zKWi0gzAqtN7jxyjoRvemVr0NIz2gHtrFqDo0v0jWOEuqGRugAIeCGots
ssMw2iHfylOZ+t8Ts4IBdEYAqeCZyNvUoKcGdII1SutI1YOBJ/hrNYlwiUqbXjRWZPpaQ+w0L8F0
V9q0QA3MoRlk4L1JUbz5XiwEZ5o/3SW1E8Aqje+DEjxwNkTbKdb5qL3w50A9kZqtqBDGHDwux5Vk
BsviwOjuVU/eHoQ112VSb2+88hVIsfYSiGM4WiOY4P/SHtZm6g1giynKYXckRVuA7fmMtTvRYaq4
0GsHiQJTiqmGghO59jZzwRXi04i6SSbxCcOnfn5w+vlJI1RbhYLg14corjzoVPYLm2EwjSm2ie5K
AUvM9QmhxeS6gj3WPaCxL604IGQjTx2x6/a28Uo4BVKa9wveuZF1XBiOEL/ue/bOWDKk6/JvUW8Y
/xSo9VsoJXkr610r9IF+29MN/uNvTx9trUErWaJZPIBVE0gsv73C3dgnEBwrkpT+BFHxE3fiYykr
Dr7gjPRs7lSZTJ4q/ShdnUSRuFikxqqCHE/HjYBJsINFYQ/aOueKRW5c6vsgirPwhuOzCtb/1uM7
RrJZ1Q8LZWMP8R2/79sNC9tIgE/5Q04OPR44IyuAv8JmiEbAICOy4XsxI0q0wPf/nmhCcIzF3uBH
Z4YNAzjmThiBAF00t5O2UhvpQ0axl1VKevBmlhIrVJwBXFqvioFKDrUVEAPSzhmpAsZMlRNDF6++
iQKQrcdg9aU9or7xwcB297XGC3BzDaN9tapkFJdRWnOOlPajcqxzkOf60TibrfT6kurH8Mb3TIAJ
gQSnUpHH+VFYbRt5L31DttCKE5UljAUH0Cw4k4Wrf0G+lRAH6+YpMUYHBjZ+T7MygZvx9+/ZHrym
7/rbkzK1ekwNKEq0OymVcxTgHZOFkcmS3cd0ql1jLRndB61IKRHwvkMNyo8HJck6Unhf8RBll6ly
BiMEOYyX8BKs8AMXsVeLhOPUv+xxyc8L6kJZ6edfhmqB/nhfZlc4HPnluMd8W+lcFne0xbxYSj+Q
ggiLTdRP3Bv4bjE3pUIUGW3O32hTsBQkLufuxZBAry28s7qrTefAFHrCI48FVllaa9+gFa7/RXYC
cUjFzHMaPNsuJtFBqqSZ2I7xJfTET7hQ25x9S60/mAtpJ5NAzaIDqowaykETqxTX/NLQHFfqi+AG
Fdh+t7JcwxP3dxMVR7lYQVa7c8Dsb1XCwRREB+axqsaDERN0NvhPjJ6Ypj8Lic0FBHBZQrIrRIl7
qxI/OHBfBEPuBLU+jUJXxxCHc6n1HGFy+GvoQAY7X2b3RjbvEB6DAYKGL41mWcQhdw+pz0raiXH5
cHbBa8bo3TwF0D2XSnH0YX8P9RShWZ27f+UBKflMPVxXCXBLEVKEHRJo0gOPtgARZQL8ujfuM/Q+
r/0Ioyqx6nbclT7pNwRqPbG+X1Ltq4dLuhCv3edJHr5uqXeBLF/ZhALYePdrG6ULh3/b74Qe1O8J
dJxENxnKmVkC5zLKfkeH/eqbTbDpEKilgBiSVc097UfWSRFoME6WeqR1yby1dQQ0ApTDH6yTmdLA
5oaAjyLxFFJP9yS+JRRpbtRWxdpKAVemYzBhELvXVRmttpn4gM3nR7dN3VT59MHwyvws4RX2TpTW
qkoxzIkkv2vnduLs50PjTwiecKl/FQhyJm5bwM/Hga2qsbQV/FZBF7S5B8Xd5Kjq5jnTHETzcCVX
kQJhtHiIB1tb1A63JBsUI8SNwvWk3tzKmR+j+nnJ6/c9pDS3zYeTRQcn64ES6kWmH5zFHH4vr9XP
oDtS9koEHe3GTcGAmwm54UE8Ns5ILB0zHUdjqJkEtFnOxbUdFQLcQLOJIImr1vwjvB00bcWEBBIt
VlU0M/vslIrIfnL+A04UJ6DiYG3SiJTZBVzTPCRTgo37xmFOy/AeE8D+AR4cXbAgsAxghNZf98bm
Uzn+SO5DRa4Y9Ahy0qsxyYdl/43RH+bwhjHtHwXJkfI8nqAv/cfYMkCDrQ+zSRk/DNiJ8cDcK0mo
OQ58w7Nd0vtZHrNJAiLRfkBP6g6HZeCxUkVhQKm+5J2zlV+u5kYC6x6sJr1S9TYQDkwDhhDbigXu
zCoWvWPveZeJNB7NlNfsseJui81/azhX8fX3qQ+QcIKFQgy111/I8ul83/2KOXeiBVxRdyU5uQx5
iYCHWGX0g+cQ6IdB4P/BU/cNPz8f7uM0lwjam7gbBKOphsmp6I06LORK54wzTck3uIUy46NRS+S0
6G00Fz06HwXQKH0R+qVb67wKuxIIEeA4WUtLYWykG4/89BXwPxqcx8eK9stnNDfrDqbkbYFh80of
FMUVB0z6/9S8HzqctnqSMc5i4O26SAYx9UMAuV6h4m/zCGawd/5Jt/TaVyxwQWPswV5rQri4KktZ
znAeo9Hlq1hz1gbS3c6CUiwSZRr9KuyKcf+n5t833hOkMqsKu7C1P6NgWRE33i27hoHikIzGDU4g
cMcu9FywUGON9Cv1GPAec3aD9GGITkYBWQ9PHGXBeeworhxbn+j6Y0Vn4k4qSJX87HS9zLU0MgLG
T/QbTaLZLbxQGZJfkcI3pl/UHOKXfX/Tggw9FoXcsIe+6JxJMWj3SSE6FU3gcpwQVsUUNb8wKrRH
jpgwPTfd9irmfYkth6Y7PyXa1QgrVG8H3dUM86Oc/1sG9BxMHHDV+3GBdgx3PhuUUYFqH0DWXzGR
wix6LrjkKGXjA1QK9b1RrsV3We+SSEePHbBVpchx6IfTN6qkCaWAOfATiBC+h5NRjpGucHi2eRgg
GOFEvvwosMBpjkc5MFux6oRlFYdOTKMyZY/gvmXM+yPFwFpGdWOgZzhBqDDCrj+IJwwGdQEoD+Fr
oq6DvXRuWlmMXsadINlBjbWaO0zCEdC0q51l4yXwMoa+njMjqPRD3oAEfVu+IREfPI8k9KeYHq0f
GlZrJvsxxngKOQGzktidO9HgwxM8Yh5X8g59wGnSgNv4+CBcHwjOrdEgrwBdbMvFL+udL+9XcLOm
cENrtg8bkCmuZt1d/oNRYlk3xz8usSa6EWUaIU4fbnsw17k45t7/tAbCyMVRzEYsOIu+HOGy9h9a
W/mPGTKg1CwwSbt+PykwkBa1/tCGR8XMtrtY9O90DtHKdwWqVnqTaUxAzOaNcVWRs4aDTEwiIk3u
J5X5CtBp3Ym3VJ7Lnr+pDEhfomUmTADve0abShZ/JEeZEFInxs71RhsGCv7+cfOJA/EHocFJgAkh
juBCsHTdXYw1aZJthfnmEyqT58ipouMaNmuvVQySWRrNJ4KKSYXagdHM8ZDfXh7ivnGkXZKlvxs+
IDQcEYmInbSDupu2Q2kGZ2a2B7zGLy3oUywhVvtvTpZ7zpzrm/PqnZYNgzqNzpraLFwaePI3E+3G
a9C8Kb+1yCDPucdAg+kiO1ahZPWmKtNB4Fhb6xqlQAhKFIyjRmTu9iamH256574UZI1PFTHi8mOo
e8URA1K4uVL8Z7brl2SmzOHScVr/NbCGZkXKZBoT5dQrhV6GtpPFFhoLM72XtT+alrPaZxEuP/jI
QSbjNu6UGuh5nsdfi5C5EKg4e54TcSsT3U2q3Nw8X9Il8sJFdekM4s0clsYhVwj+0XWZR0ni3G2W
9WdAX/o6YMYrqDLFbg6M0t8mUnn1Jmd/Ha/1+PJ0nfJBANaJIk9KQiTGMMuDHCz5jXnJisTY2sQz
rigBabIgm6BBLaJJKPiUGF4ejDqSsSLGIB6czm5q0v5GaUzGx0L0qr9bghGBemiDYjOHBqCDcaSA
CFLqhey37EKzjDoCNHRwSN1KzhAHCn0LmfeQmTIpaFR8jl6dEmIWtJHdsIwMJ3dnKdbWgCjBvhZf
Q5ErY4axfpaBqPHPHehVBxAEsLngRm/u73I1Y0eTCMgf4zEyD+EmTXK1Cc8KWp2hV3feCp1xouZc
YCqMzWcKM31xgOWoHp4rmlCWqLP8mGjw4/aYK+bCbA2E7WFJ/IVEskGm61q8Y250Kz109qRMczfN
Idq/BjBgtSET2DYktXEvB8RxamTCK1U5a+WGoBct+SxrTjJkCUmVQwZ9+wDbVfxt6HyjvWV2PPUZ
iw4E3Dk6aR6KeWlYSEtHbvnrD13Qjz6BAl4BcOOMpbFMTfXn84pWIts7eQ/JW9fMSkWIdfo2BEU7
XmZpLqgP76YLKTM/AiVblnSN1rQMs1VlMhsPpzNvzxox3HQrhmpLu/3A0PWpliJKyx9LCQrV7SWh
rwAkWFYPC2ef8MK4UB3O2LuCNicN2GF56J7YTaM/de4+5OZDjpMlL+R0H4HhZNTsC5SPqcf1zCku
gptd2ggNsXh2r7lqDnfzy+4j2jICyrx7AHUOvGyig3ZCQQ4lSyUnjRPw0Q7MpfE6B7M3+WlmHlGg
2EZn38V3KIxtWI0iWVrpZpyb5C9nxb7hSSS6bwdiEQOb3c1q8DJKrb4tf0+rsazjQyMTGSyfy5ng
T3ojFQXpkklZbjIX6aP/Ik/yZ6EZ95pet33HYGbJInwVtP9plzqxbeJizTSoMh0jFAoFGJY8bwFy
d0BeRT558tjb+j27zusB6BduNfhm8p3aBLyjTCO5MHky9PXK/2f4tSW/de41FSQksVkkXkZurkp0
3LAVf80EOZYtsFb0F6x8BlN+fys9B6aFY/n/wsxyOsMeSZQ0wkezLSM4LujEtf9qzDs7sMnfG+jk
EB8Qty/YoCHuy7sOskNTUMl2gqDjRZ+Usqvxphp7uEoLVnAdpur7mnGL29/06L4O6/gvkSvC7lAP
bUf775HknGVFUCr4gduyh7N4xajT5IYquU6qfVSTy54Fx/2MRdmIt4zi34MJOKYnbxEd72lBiQUb
FamLkyb1AoKinEL90P/j/kJhUTVPMy1FoPZAZPwfwc9PP1ke58ysXCuFj9frkZHzebk+ORhq1y9l
a8G/xehNE4Kp1CwQWxYHlWXLjwiR4H6gq4DjWnS6vzj/j0FxUQ/Be4w//n7NdLf/A3fynEVvXfo5
/OC6ynWPD/tOTCNHfF3rw8OthZKz8brS7UFbNZWxkGWVxWL1IeKRyc/DUMlC6utrIcvUJ/NmU8zD
i7g0ZrkVP7CsvEBqo5OSLuhea1ostYxjyTOtbORGXAfihczuAzYjyN91gEJc4E5a/HmIzTxZiKxb
iNBmoc9+bllEVbFC7SZmuv4/TTU3UbtOsiUo2Vp+ZalZH3WNQcfR3x/586SRlsHFw2RtxSACHn3b
QlERCPZq94xMQxQ1KxXxwcAgFVeNm9BrUxn8jf7vyzKyiSA8DPOTgYHTOHq4okrlMg3jVbYl78k+
eUgN3JaqmVcwfdWBlhDaEpzYRrAoyuJn1KwvW/fqBt+tVVKIIrH7CI/oRsqEbnZrwOTF3LZhU3bg
Xa7R/r4wtYLC5dPCZ/9W2vfrCAEs2b+yO/z84kQ7U1xgdSYmERMQzVZt0P8D0/+43tdUNsw1usI3
rVHU/4lLSWTQK5U46uNuzHQhEVWtfrOKKDTtVxpxK1MdrFDlxtr1QXtcKWLy/gsKltKy9dd8VOOt
TOJGK2B10KddXxiUnrSQZMgIyAyj8C/Pf6QpGn+wQxKTURpg4hu/+o8URUaFD6GvWe4M2bHPjx++
oCpU7YmOkaDtdey16HXhpH5Ov8hgwQc/sOrUQWcCbecbCuDCSkWtMo7K04jD+ZU/PXZ/pGHie22X
od9+VPxzdsj2mq+1jyXL+DDK+nzq/jrAs/0cKVZyCh1qJTPPIVMe6bdOh17euT/DkZo8aRHi+8wM
CNZODEHmWrCtzS+0o+OtMRPB98riPERM+qlXh/heNpAfbD5Y4MGSlSiY3sW7z3HcYVYXJD5XKnfo
KIxL2LaNmfOwGFp1jwxTr5nGsB5JV/63GRrHF09VhM/VjkLq5pcjcjLQeYs+MKKa4M3ZGgYQk5UQ
v4K77rmwvOGz+0YTwGAct5Rzd47etEXsqerC7eHDo/ancxCdfRaX2+aNHXP1F3UxWH7iVu4BM15B
pXetc1fJif5GnSRNyIL++U0WBBN1G8s7TfhG4B0HSxDDzBrcRnfniMU2uLhjamUMx73zfCUrMOlJ
5HclMsGY07sukJd4yEs0mZgnsMsS1uS8gcISe0zKYRLEQ75SakALW0WuQaVfszimpwaKq79yUoTI
PyK/6CuVhIcv+Q4VyZTp8+CIIKNivSlLH1WUZ7GSnmiAjTpoc5uH5A19EPVdORdwtD7LQOxgXSEd
zVkvVlUf7jYeNCg3JWFlHpLbsq+wPHxe9GHIOEdgw83iWdNyIENFfPNMC4NCjfkDRrKirKRHTHTy
2TumFjbHNqW1Uuc2YiYYtrTSDIo+dg3ce4T/d5S4hjSdanq0IU0kl6OebvTweNkaOsvBmeRKwj38
pG5baDzzgDBIMJrVDlEqBYrOp6sWk0NR2R2qGZ5ZpxlEh4e4jchKkvlVRfRSylP832+MT08SUdBZ
CKVezz8XiN09rWJ9Nsfhl/50yX53xaOgwVaw7L9gdwxDldTHHhIjUgdZaEik0/NvznUnEH052bpN
ti70zbOyH1T4IdyaHbmccoMKDbpTDK9qXlaDO/jzuP4svfEtVHze2J/coMPrImamSsYMMMojj4Ha
H01G3hVf5lxRiPoAdMxeU7jfrebOdie1AXusw4KoiwI2ieMVLBkT7+VMCsqcG0lF1vnsazOddt7Y
l2tstJceP0EaH/TUr1iaGnonOYN66d7Mrfn8yfj7NdtUPfphqc3Hs96ZIP7CWtacLWpnEc9S6Wrf
msP0TKueU0C6HXZa166qClkgDDEDN5pO8dEmpMlTceSxSY1ztLs3RsW9Xbr4kIT+4nNZ7MWasiNi
g2WBghg2LMR/4CKgMolnsd06EJ3dCP7/KXWIVB508KMysgPd3jKQ07dyP5YOweClz2v3v6Hte/qn
C7irUSYHpS9TYIF7BCBRdRVsaMlZJ7vFxDjNK67o5WMA7TISqGKece8PfPnYhSRqU2HKGE1UtK13
z3iHiQ6xEKiDVHFxsfMieuOieE7UG5a/noVcDegJr19AEkL0fgeVY80v7z5j2qrrkiPItkfsOLBJ
BwWhRvMPZoVOHYchJqn+BVNUi0TFXJX3uBm87ZaUEPE0ElfqeiAREaPdUr5n2bNgI14XGqyJ7Xak
s0P+KAmrX4IOn407lK5esWZR9MQDUH4l+EWNkvzEzW/0D4ajTjENsGGiwB/XdaRRzRJr3iImVrP8
fFK+2Uz+pdvZK18kX8FXsIBvuOUGKJIWn7Ajh/VPk5/6aqE+I5m1SSNDq4cGsQxSghsEzrC7LUwq
Wt/oa+yoApDk9xEO3Sb56EAXQzdKiQnwsN+kE46HLmtFDxg3/vIvQ4+p5TbvIftBX/YsyOeVzw8J
OViVVI7UO1lSWfunUQUbeEUlmX5p5/quuJG1dAVQVrkEu9z8kin5JnZUmIyBGD+9+AdH/GyD36/N
HN/e2d50d8jyVE3sRn3pA9Yz3iOlAfpf3tAbhbZmx7yYqrHpO8srEPrpVc6xa9mgKq+l0rmsVoQj
uiWewawwrr4dcAW8tQD00B1hjV/mvbkWcM2q3x2ocIR+qY8MZ9DB+VHPteURCR+WA/70R8ydkNZo
vc0CHgwZTPKPvQFw2hPC4Nh5dXkQPsnG1TeeFTU/Hq+Ol/rlaQ4VUHdYBB8ygbdU0m/WP+gD2ZHY
47/ZAAalCMZu7hspUKgHZTK6wmRKyITNWisZZybAUd41AGRvZzWbrs1Y4/D1wjoDvWfWFXMmDYJ1
ISeAS0Bp8zvnfayjr5EUT1O7EziWab7MLqjBx7qPzBme4z+M3cvE2e6Qjz1Ubu4nkmH23iTe00zw
Z/+oNt1oCtd33iV+6Ew5Lxzi5z8ALlrvO3yKpAvs1e4dgYXcvF3d+np8XyIZn6soOSlB2SA34PCw
j7nxpogVTC+aqziSTZk9dIwv/DnKLOV5efqB1MVCTQ+MteZ8yNGS3A36LZ8F5fhjb/k6fvq/ITlB
PHYevKJRm5cv1ynhoSzKezBFHnEl6uF9Dp6kRCLUeEYmsR0dHRkmnTOenZoLMsa/g4J9uuV1c955
zkINNE1DHS+xzqR1Ke1a/t8akucTe6jE5WpdocnjzNCFaptMU+TPp0u8PUJU8yhued/4WW1MNOgc
Zwozj/DDYXU1X9iMaeH1hSRjOupfxt2cHfSHR2KFwwN5v7sRZ3b4a532McBnZW9KhEk7ecVox2MG
SQ7BH+XgAGbecqNre03ymP5BJBfvNzEvcMJqgY36fOzdnIzm/Cfn8NZ9lboPc7WaHOnMfLDfm0pG
azXmDpSQ/oRKI5LiL5NvoCFwTTJfmeLAPZE5gKcKQfsglAQZDnwpbulgDtFn9V0+YTyhsZVEWaHO
PckO1xuoCpljdjhshvtoXsyrnizgoRx6JYD/IUzDCL+VefNJitKPr4t4ariwBdaQmWaDOL3opOU2
4frznWi/Duu0aBpyhqOlWQ+CvxZTF/W7cV+y37DdBmc8727BoFzHcMpemIQSuEwsiyzVvbE7d98F
Y0J11ky0Vq3z4EmTnemmzaErK5H1KrQIdn22zt7ZcxQ1T3GUPfhX7bcMSopTrN8yAgzL/LvhqQy5
OsyJozrrH119fsn5sM0Vi/YkrMK2+JzYFAIcmsoFGuFREPxXmaDiVg5XkSeieGfymNo04iybWfqf
uQOcng+zIc3emVtvSonMJ8HnACx3JhxL5/AmyEnzlvbDA85DwPgEvZYf9R0OGK3JyvoGjxtWCWRl
+MIvmle5JYaItSL0qlpc8sNWS0G0e2RH6P1vBVi1sHORa1dLi77RHqrTD8v+Fy7Kpv5IifZIyvQU
qS5fniUf32nJJGTrRlZaz2Y8I5mcLKC8hfJDb/Y2WhAVnCNvZQn86ld9OnU+qm7g5BfTCFNgXHBm
CH0mji9t3jjWwyRs2L1177U2vQ68le6eOPyMkoZXxG+GkvNaKgWFUbDqqMuAh9R9htGJxjWjA+8C
4ktiu/sHzomKIaOT3fU3+MClP4E9by4YJbreH2iXsHx7R1HEx97wu3QL3c++HRXbTJQXPDpS1P2l
tnn7qVPVo2ropXiFo1ux2UG5doFCAbrlAPWT5MLwPeW8ScgoC4MCdlLTUWz5WxgQ2VCU5nTERzS6
YcZk0zaPz7CuvXf3Bpt6+gdNRG0HqFVxOMZF+T5fdkpzI2OvQOAeH3J8QyfqLviR0UKa0cz4AzTf
gNsuec4R3943/JOEsdufqFuK3bY5iTwBla4aDhMbyIAwRGtHXoiGOCs0Dv086JZu5AgRScSQqfcB
AWcSHxAFp5Bm+MnPnh828reo236c2BfpNk6h6d0ZqPEf2Idqt8Hdrj6qYbNPVt9he5Isej2x2w5Z
pFW9LMBm5JXFGMkQL75IlUdCr7WSYmfcI1/BEkaFuqWfQZ5qXXPiBEg5HEumzawEDW4SWm1h0Uj0
AE73AlsOReKCTtSIqJ7w9LxGLbkw7VnnPdcaVXGjXRjAyKZB/bc3FZr8mj7VJYgb52kKEvbG2+Ir
1JFThSaPMk6KxboRVRoPq1MyAO6pF027KNwF2+eaH8r4RBvQ8niY2/x6V66l9fy5mkzPy7z/Q70s
AwEw0LSQkvwje7bH3V3s8d6gx3JaStFtlqFfXux1YPSBZeUsJAdH/777CaYbhApUl7Ir+Lzc9RDh
F2FmlC2jpGfAwMIhmRLdjEyMZXFdZRK+6tJT33tRfZWW11zFm0devsJqUGlyIhXIlooaaobZb1iJ
Gw6i2vUy2A/Ywr/hnsPvHGox3vnZ6tKDyqfcPaOBpkMXzN2AJKpWIrpXrvCr7TK2UGnXLnFQLLB6
Ksa7gGYQnx6CT6jthOVwDLzRgOVKyi8kF+BqBZSqyXAWi7h1WfR4lwnDsy3gg1C0ru4uJTnJqckH
YbB0EfuiZli8JBzlNLwEioEL6vYnssyY9/eTACimMQTDYvLM1nUw7CZLna0IU1HxZaPDkUQuIcUz
XqL6pa/nKJ38Mdmyo/vE7VO1P+dpXlG0l0YffYR2bPewPP6LpfMib9+gKLkEZWgNCzaIRNR8j1VX
jJwPDvnMAH6qTdr9s2TV+kYSPAoK0WQQB1PzsKaqzJKXW0xm5SekM5mBWlwje07nLDhGoGkTIOuu
dJpKxi0JCseumXAd9lD+QIDWk7kau+Za6xBiiMwuG+zLF3KWfZtTntTYC2uj5sVSwfEhgP2liPrb
YSE60z42wDiHn253LcaAiR5ztr8Dhx4504qUUGrpn2Ph8z1m0OO85tJ1tRu48x8e/oziWkui65qz
6gOp9Ve5AMgLMmj5b2G976fWb/4URm/FfXebN47YufyN2UGHw850liF4S1gvOAPY+eu31x+Zj+6n
QSaMzLevn7nbF2XTqHPDPgR9NwO7FQX7WKCdGgZINIJw2/Ddhl3MX3GzfvO8pQKxaOimcT3+IMg0
0JhKkvoDeNSFdEm4rxjx8G43fiLbOqB6yqK8ffT5uTBipkPi8LEN7PY6iEidyA+o4kgcQYGNFoG8
hDUO6935OLhyvm3cqS877NcJD1HzgVcBnyQu6v0nElrWlZ2URzq2w28ZbXKlkvgRQDEHzB21brWE
u3oWmb6iETk5OfP0NioerX8nk1EVgS8vJ4E0w8teHsbMVePWmypqazT5DHOPlzk/X4HJejQ6TVC1
ZdG+cnFVrNYZAiyJOglv8GFkX3rbmpUXoDCMPogmBb4wal1ottLOK3ZsaxwLBNIO6SnsG1CKw2sY
KuwLyBDP8RwxHUq/EHEBfVBsPWgphc6SBRiFKNnHB/EMo5uMLyhqoAAnMNnkfS+JC+mCBbqcV3pp
7XNRf6CFm/coKU8f0IA+DDFlTXZEWEcRFHj6qxQMtfKgUAh4vbOmWAxJkmzG2HWvzNn1GnRFM91z
z8BjrDk3cI0lLxSeD6HkMfS3gVv+TCgFuQOK1qSnEPsXr3/jHbk7Z+2OSklx9ieJeq3omw52YErF
UkkGO/o0/wCkonp/+9x5/uAOANSx/gdw0ckXmnu1Vk40WtG7MzOkLyRwsEpaYNkzdkeXflR9QexN
7u1y9OyRnAPM/QUE5kjN4nYDmV0npMBOLisSjD5xvibI7o6sP27bTjEEXMOOWXDwN5ioApW4p7B9
g4kNNcVI6onOC8yqiGw1Q7+vYY4uXNkI6gRQDx0gF04J2vCy58K2aU3ISxS75HfiNornHr5vOsGj
DHv5bq2yk15XmCbEXEYWmXluqRAEXksZ85itCZjLwSHyLStelgEd0whTMLr+iWgUEG5YOHKOB4R2
y1PcXq85SmsxRsSdgSvIbiSE4sTfxFnCgzkOyXUj8JzNL1BKA7INofC/ybRtmnOl4hYGaN8PyJW+
Vp7xmWEBEgROeWMapZzyaxgA6C78z6t8qMdICmKzNhU7OE+y9IVpD2qTrtidZZ+h4z2xWRUzz/lN
SMjAyXkiUr1LxYEyGqyjoW+8isXDvNeo5sQIkpDDJ+9Ly4suQk18Xwy/MKkBrgdCWqfnaAwZyTxq
yc1kM6GO7L1luZySlM2FD09lNOwAmOoDis6prQMhPrJzOVT1b63PcKkhl/16OMVRB12/wZfCgHgL
N0GEPXJuiKfe53n/h8JMeQw4ISqfM772869uYJ1R+QuLlk2v52hWV8f3dzruu2U5HBAtzOOr/Rnx
MdhdcBq9MSx77pWx6t/Be2stPKvbLlS5TfyxiOUDMfjFwqMGUYNWUW+QuiVgEQUrVAyF37y6sMJX
PqHERtI9X8WOPki1Wgg1NsGYEdHLCgXNuyiNvvUmyyJZQdKvH5zlu8geeWsHhpCbhmT8zqYl0sHM
zM3HFKTo9555Iver8oe3lY5V9/jA72g15HdkUlDyKEc4VrYCHVRgyAZPx2Gr91huokayz1+3m9N4
V0ezaSpPVxCX+kZYnycFmT3sYvQkwmkHHKI0EORj++gkQEeO2OHBHoEMYaCJtFwe+aMJdFBPDbSV
yxml1a7D4E3xyqd9e/iM+X1Y6d5lMqJKgMztEAVXYQ91Jkaxlk2D/BwUOqTU0ibPJn2xLDBr8z0/
aT0zZT3X05VfEXkSeoGfvuuzZ6HSMRijPBSn2UMgbb1yOSAVbC36gnnntxysabGerPwuw6uOqDcB
uL6ylehDwt9ebjh1E7l8doDe6T9H+28FNCykOUPap/husim9q0bMGnLOzrjcmxY0/9m2tZQa38/7
nK75IHNCQNGmEvI1tSsA+JCWkQhcXMfzi8QOvVIRYzqd7IFDCW17ntdPPoEEUFwQVNYqvA4xCCJq
r4srZLjgj14vUFqP4C4hnUPLSbGGkbwUAlqahQjiGDXfN33ZRWxZoPpcfjzBOHPdxTggs6Y5ATgO
sk8c8Gngi+BvKp9GS/ykC5cdnjF/nEj9pRmnnb4cyEkDXPDg0TeYKyWzSLY5Td5QPWOslYVUUXs8
2F3T/xQp509DUAhh4TVTPadB1SJ1wQytRMNvlPPGso60YM4uVj8SoHhp4Ojr20JWaiHX6z2N3vy3
X2w7nsJEeLDvvYC52fOM4YR/jR922gyeX+8743nnaKNgbVrripF+mHPjk47sORADNHCOxPiiu0aa
Y9I2nBtffMIW3IdkMlaiEljJzf8jLqfDSbmhBcsMcMYRE8PQOdcedLHsXHwZcGU1rk5MUFfbfLRK
9CG2PS44N3tj8kDE4mIJQKbuOLY2hnhOSgHxcsm98bq2EG6F8ban1wqhoin1d9vF3fQb8HT4jWwf
qmqO43ABWhp9RFuK9Iw4ngGaRRYnpOXHZt4+UndoSQ5PKHc5qek1SKay1rNjRXt+XZifLN4hnQfk
tIJ/Fl6Kv8OKNDSpKC8MAecab1Z+l5u5wVsz4xZXg7sg1d9UlanIl9mCF+0wt3A8LEBoNiiqTaca
ke+g/I3OYx9D+3WZuNrSLyw3wlcEgzx8upsexn7KQI3johem6/YLDpo7U5I7L7V+/52PGnhKD5Vu
du+Gb/VARlbBq/Ht/YHtgPAKIRPJPdFQQdROW1I+HHIhoP2YICJqehjVq9gUXbzXlgvHe19HWcs0
vDcRCq1vXpaUzRi1xB7zeMUc9Mjs/olkH/xaM54Ddy6Ub1uRarP9uETvVLhzfJQOaR+cQqLGMGbo
R7gMCXj+J6fQmElofDfbyuciZpNA4Y6elveDF+e8IgK5x5MkcnZMIifWuIejFRJJppJtU92A29kz
2TvqT90IlOhY65wXJP8RG3NY0N/qiLhf8dWICi6OUQGcCVnrPh6rJ3zu7hE+2yaioHmlvCmx9jwz
9DUTSRLPT96dtc5GtO7x2cOXTGxotJS3u4/nZvrLkv9jEpxGCK292V+NaHhveDj0GJnuLpaUFxir
pUUjmYvLbK8jLBe1mjS3AXDNNHlYYqfxQ9DJ6EkMzZRKlvV2/R0/U0pj1cRfPc/XTmHWr2RYrSzJ
Bn2YXftnHeMC+V8Sd05ySHyqO7YaxX4ReeUgDZuaKuLuPejbVfSEZs+s/zH6H5dOpZXbLmyZPR2F
E+qWXWjZc8Sq2NeMNNT0c753aSO+U5hdaNFbnHDzoAkVGGG50ocZx1VHqHz8oiYOJN99OBO3aTY+
rUG5Z7iz/7i4++sL+uPVsVFYdqGaIENhs1BVadIn19JVdWV/P8TqMpTfl8vvcMyb3IY4qsL2ZF0l
2H3l4/oU82gsBiVI4tPKcSVqx7Q3UCdSEt8g5a6qPt7VERGjGgCqzn4ia2kLg0/WAJyJM9PYPFeg
jgFTSAgN58/IqcpWUfSz+18BXCeMLFuZfluPeqLPsYQcKwj6eInF/a8JzSSOC+wr8eSHk/m9tEhm
12n8ET8jDxqsBurJ9rptw+/RFnOWLHysUhUi/5V7+t0Y1GblT8fmbWq7lik0diF5WFybnKoWAf0s
XVu40I3+wEWfa3avx0sPkaWXhhw4EkU8Q+6MbM+JwDvjPemadUkUWxRZob5BMs4d7s03lZZ0Zlps
KjMPQT8rHIwXHrOb2y71Kz93J3EyKiB5j8QuK8I+Vd2AU29XEuAxkbRJkOdZM4oF9SsAN3FrGTJ1
Doi+nyCjzak/0Ydgd6cJ4uIo0nk5xgGeIs1SzQLw+Hw6B1CehyhocJo1IVagSbxlembjmQulqylU
XxRDqNSe4pDIXDpgXzmMuYkVnClvwtRGKunC63TSzlaL1UgUBmXeHCVzpyYAJTSHMfiBoRNrotZY
ZOyOeRRCtQQwpnwUUUk0qmmK3DNnVKuXjheBb7Kfh6UcYeHU9hUXPa8jYIgBllG2xDdy9Oc42Gwk
CEjbWGFRMxuavmdHT2iJa+QE02/nljcaXfBRpwuj7th9Be188ZY/VWiZAj0WBIuE0LnhMrexqU90
CmL+pfGusVN2mNcAAd4BmflIp7deijMCKF9SOHDJkNUBof/jspryF56n1+Pv2r5wVO4SXnbNzPNk
3m/TgYDzlNO6U3ZDAa1JUjrlr3kCAsGwluKRz4cPO2mHkyH0gPPE8jibpnAgd1+Fc0VOc8IOUCsb
EnBSVK1RYYRYWOSO5qx+JpEfUHeyLbbK8arvkS2gM/NJPDLWaWY/6T9qpEgeQs7xUhZ6QVw5WHDi
3ARgetn9AxaVrbksyMlJfNcK6T0Lw9+lGP20yUwSafzK6aBfJo0ED3CaFgqTGPPGKAebuI146G+4
jdsOYh2kZ8aOrjjEbFa/Ky0y4VWU/0+oIOR9inhZ2zzbGu1fu9vB8jyMoNlzU28jkQrXjU/GeQBL
bb81cgS7zy5wFMdVX0iZLKP6nP5bxXcaJAAnX1AUYxRuXhd4z/vfDXnNognKNAM9CGRwGBpaaT8P
ZHnGSuLSPcuEKDXcsdDf/K3fmSQ9slln+Eazu+h4ksbNy4YhvzjQUgutaRKUPHbHVELJlvXXV2uz
kYYXZjm6Tgs+8gqEsCdHlMrCblg7SPaFfUUOUK5Izbj2PfHJFL5yKwWmsgfplGabKVJxlVWQOSIu
7yGGoTIx1mpmG7xRFz+cAZ7H3lUFmFpXvFysvCWm/ad9oLmtsWc3IehbOcnMt6tV1kQ6RW9wYmMP
MHmeN5CCVLAId71kGVbod9Zl+LsEMXZCdAL39HCfpsI//WpOoJxYZ+PV/eB3S+JavxNy7B5Miibc
Wvazxj/IpukcbuhdxgR0ncZzjU3OnrLKGdwIdVDCCHQRvnsadDm3Qd1+vQph/wfh4Pq3SPfSKGnr
zMXe4Gr/HnKJIDvu8NJLKllncOB7wx+BHGo0dStlXXYmTsmhEuvEHHQT4HOCg+ALAo7flPBR4aQ6
cnkFJM5ZjP28IdCfHMH5oldlSYuPZeSOpTp+KuScydlJ9doSwgiO+5lu71l1CqDnvFoTJVpy/HJf
12wH6hvNbjq8ELG9YclzcAx8aK18OiaOMwucLkaUZn78/Ae1PNWfpC8jHDjj+9YZxcxKKPF4aD/t
Ntbbqgjn7HttjvNY9cAh3AHqKBIIAQdLbfyiMlCKb9GEt6H7v9HkIcgXskE61H0Lh04X29vA+rbe
J7p1lD9Po1koZEh1LoQfTK9SZoCVHVzFq5qOh2m7cJMsONRk3+Ed7pGLCX3PwPZIjIjv0g0ngEi/
DxMc3Ng1soNfp9MmwjebfnmsJsSBAvqPSRmGqu04rmB1wWhnco95ZqxALpvzgJQYPr+FMv7dxLTc
P6EjRM8JlVsrRRS0IK3AXOjf3/NVVKt2hJkwLx8AMz1ez+r6GlceIMZ4MQuPSeTPGJyklG80hyu+
8Nxv8nEJCr3p3SdTq5CS6oqxHXA478RxZBiVgLP/tcwFav9gDQv1fsH8VqF2bal6ZhfIIlPhZcud
Sg2SMrY4JCYUzv/bT84ZGM80Kr1ZusClKlpfI9VCca6HnOzeCiM9Xw6b8J3UAaGgeQ0OJn1CE4n1
iAeaS5eB11Cs5qb/XeWUqqk4S4AfAtpImofYs+VhNrRvXCpbuFf/15Pe5GvkQmT1phcl6EhQ3r7s
rKlHs/cTWS5X3OzGT39R02W2J0lf2cvmGis/guTTiYsmN5TUDWjhh7vR2Zd2zFC3lr86Fe66e5SV
llLyL/gUnvy0YSA6cFZRTbmDoGB5XrVkH41/Cxoxx1JWblHWiH46lbedqwXWmrXWOWX52wsIU/yk
OxrmOtQjflbbtmeqckMJg5v3DbVV92mnh5RIuhtcFr6M+M7o+WF3QG8qFyOlHBfKYj2M7RR+kW3t
FCvUUNVWDqHLusgPT7aLVOYgm+NH473TsFq/o/o6CU/afCsnqGPJJARuTe8g85k3tg3JHnyiq2ku
yxJ0RHy2gi7kSZDuk9BsrrCRMNMggOUXeZgXVMYOtXA0asgCzrUEY/j8YChizZ6gj7ePe11lHDDZ
M1W2W/OP/phDD62pMyRfj8SY+yVWRo0hHGsGhjQ48BnTbUKQnvSuIDUZ+gvJpTqIq8oFSz3w9Wab
J0uduZHP2i/XmLSmZxSNmYGW78cORtTaPuCtbIF7qyjsHqADi++/7uapQBOPYB9PRrWTqeAp4W8y
CDPUUWGXhJXKnC0I87GlQFqrc9UmUTE45D9IgQeowygu6WGiUkkmYmWBNHDEpmAHZ1Q0hExgYG5W
vap3KhMrHqa4uqpI111zCXHLrQl8t0wTcE5CVlyXDDxdQR8YtNGvldTrXkGhwOw2fKv0+kFxCGv5
FKp9H5Vfy3okCwua9CCmZs+yUbzdLEAKSyW2Ahq6v4JEKVsN3K9BkJqGTGH1poVHkleN1hTwOKXG
SvjCYItURzyZGORqTY4s4fMUmuYpJB9zk42qSfySh3wbE1ntHZ8FIVPXTMCJYv4bBUFpuNOdk78A
juNdMzCg82RaDa2XyGI1n/9ASgEC3y5QX23oCsj91v5cVNC8rDmYMqyBhB0Xbdqq84UFpjI3aGYH
6puxSDryUJqMc/uahKHX8q8gPXEj5YijqN3x6Ezsgl3BfHcS45HGcPREWuZC2vuxoJwIeXxb37wY
lwml4/jb8pdqkzYWZP5hNaFsnTzPXZPVBhMj1hLSlBTeg3sK/Pra1MouEHQOJYqDYRbBUiKKE/78
9sAPaYhp1ZOiA4CJ4uHjE0V4Vt37An7Rk5EB+tsy3HBV3LpVMbsPNGp0o2GJcgUiRkvgslDuudzq
iEO6c89veUkS11uwqMg0VG+zPMSQ7/cvVvRatQegsw6rerqOrr2/E0O97JriONTg4Yd0p4Lt/3g3
bCs6SyEi3kvgEMvJNA5NkwrGCDq60mHZeEvHq401lqv4y6KMruwz09FoXPKzJawcwQw2ACN6qmPY
4bcm6y+0O8XnUUMEbzGPTKaD7zSD7gwegBrFLovA3HKoVV13G/pGWfsgzqssWXnHC7sSkefjxx+A
//qnVwkkOmYv9aRyHtLZtTh2ElU0/cwFn7MydhbFXgMrg+HF9YVXZ4D8PrTwtmMsUPWmFYs53X6d
yqP4LWmRv/lALU8Lfl2XDJxHWjXVaSDEHwqW8sa3KRZ96NpKJJ43wndsnDlw0Tr0Gq1heKOCkT7D
+Q44xJ+0TG4RBgLVEoUstuZCUAaIauufyJD12Q5CjrxundpWSOxGMb+ZViBwCBS4M3i01D6ceGko
D23PweebdWFkanDJJ47r4pYStpIF2Iw5zOaDc3C3pHQjbvQGL11M/gb+h34xRcG+8UraKH0Vd7il
9UGmllyKVEE3AG4ZKBJGzXAtpx8WdE5QG+howAhH3P8G+pTPGeDiU7kUlFxmxr2dErnJhCWVTDjo
35cP0NHRsKaB2/Ok2G+XNMJze8Eg+aNs8f0If+xljntwFMHVeN04Jfmt2JPE6pVb23OFGetrpdbj
ZX6dX9hyHI5vpZ2gbDVS/f+dqAC50urGhn+A+O+ZrCckgYZuaCt+zcbgOVDklgKxokhm9v5MNRmB
0rmcDrVmWddpZH4KYdpBh55xcj+vxD+32nolHQAoNrOIaTWiJrlnuSya5kPv2VbgTvqrzVMQcj/m
pAJayayLR/jiHuDhSoGs1HnQbbnnwXrEskAbcdgdKUx2oE3fKhgbqVRj9dmOZdJNtbvrZGmHKLw6
bRO0nSRHRs3lycJzqzfLk7uG5EKLUsV0ddfpZQXglRrRZbBOPqFKF2CEQpbA5WIbrLJaURaBbqr7
0FByyOnX66Stn92yX50HyZsTvS/SHxs4RQYiec/Qu5iBMh6d6UhTZEAV4dUQefM74G4zXOuLhZrb
ChTX772VG/TMJ1f+DrDL71HstISWITQQ4nm7sjTzokXt58aWGxEKtRB/G2AVBUEd+pJ00/EbkehM
leMJzTMqxCRTP7OHkKobaWJB1Nfoceo5h20ZVKDQrx3hKAWrQGtMbgZxa9cwz7I75ND33vC5e3yQ
vRZZQu5mWEKXPEp36v91NxIdbng3hMSPJLLqA/UxGPvIn80zxjZq6sHgU7VkZP7ljHkRgR/iL8Jr
DbVTTCQrqbof/HxeWdbCNi+vyaalWdz8EPq95nWNXgmnpXT032PgHY0XRBZjjekNEAq+mDALH8Fv
q0IkFCFQpo9Pv+nbEe/wHskcrHhID10Hb/gX28z5MPsV7mSfL/FvdCKzXTKXAf8TaMFLh5EwS+Ne
kJ6Tqc1ckZOLwr4eq2/B/f1q5Cj2B0CBo0AeOPmX0QQuHXEzqsf9O7p7AKcqEYlPfzMGGwouYCbh
CnyweytLa20utwchtAKectf+RFKtid9qlT1OmdH8D66BaPMBYdl1O0uX0xqPyYaPumxtZTf23Mm4
Xn/7Te9CYn5wedcxxvFN5Ylyl14zeIdSCUo1RwGQtPRqD0P7mEaRPZ4ymiXcCa+UPotgp+WMyUf+
lq1igCIkZE/fBeCfKDSOjlaGY6gWVhm8P17WIVeSF7PABo8I8Nt2n69B8CYLKostkzST4eNVEaAU
cQwXpvD/X1Hq/33RkhOJr6PolpHRlnCYv15FCrm+7g7kNDbip0x14ZvC+UNvH57b+dMeosdHGbAs
m/7+J/BPBl7I/h7qOmQtmq6zpACDas0DLPOCYamgkZyHrWbofYA2E8ioVUACmSDfiznvoD8VH2HX
tyaX/lvRnmrInwu5Oqp5IqztmZyYU5ShJ0lG5yh0Ybc/yHluTx+9Za9cxFgm6UkVopcn5rmySpxB
mZdP/1lxLW7BpF11dbTTcuhnbMX/ThSiQhAaLWQGZ7GIT4EAg6JyVIGyxep5r4rlV95Mhw7EQd+B
SRs6VChPC7Tg5KIBXZSX4XaTM8eoiK0ugQ+lcGKRCPwJH8eI4fSLHKYq4PJNARiOVYqmdlCgH4cy
cZvm2/y0V7Sw4F9syKVrkKutoD9Xsat/HLyajUoO5o0SUEaB3X2vozrsl3BUDFU1cjZQEIhX+gBN
2gE0DDi0TDuqQd7/fPQRnBGhPzTe7BjH0Hgmx8lhFHpjsyFFL2op9pHV0724ovzQv1NyssMgg6GU
WS7UnliNn8YV1LrBBZJMoxa5an/RqAAyUdEoTXQIOlxc9MbiJDldMvMwyK2BEOSTHOPJ+5hfA0Tc
g+rVLIYL9YsCGxZQwRZCnsUWK8VZdmwF1cvVMzc5nM6luSPtlAfSpn99QHUOH6689Ysr12W5agdq
/r8Ft4nOQMthO0kJkuMbXUQm6AJHHvL7+o4cQa9S/Ow2SCJxF3KMfQXD4jRk0z/lEFwUs2l6mE0W
zMYSqAuOObMk4cXQfmTYh2hs4w1XtZZ7sE53eDSDjsJEysMLWNRO+2dygqljtM1qudCk33uJ4czc
vM+vKmh4j+cQQGegdnjIHYe0fd2LZ4Dd/5yhzjb8fHbCZfdGQqFhoMWwZ0q05rgItLWUsH6nNfHe
tL0YOgMoPWg3otUuqYPNS4+xG/P+BwNeXy8BwN3tpIgY2rf/FyC9p4Ms4QgqVcdVot9DA8qXuyyI
4Ci1v5pWSchm2bzD25f0xmtlUk8iYRNCezHhBiukT5nKfniYGMlcKq8cRgJltYFujJTNyD4VjDF5
QJZAJT/VYmEzXlj/pRWkkyttQG0s8qrxpaJ291MdDS4zEfgMMUzglv4I436IZrS8BHlKQKKGNpBN
Rr8XuvbO8tD04dYgjZ8qPx008cON0hpDmPCDXxYSMUBrjF17VTPlgSAB7m0m8dCdeNFTQIBNv738
zSy4nqY3Gd8U/foXOr98INX4DWGFjg7Z4sXczX0SYbossOxjHRPxjnQCY50dQvzRGp87VBKlCmG2
Nd0K+xmJYeMVS6Dp4UoxcvXxi5uy8Gm2qaBbfXXxgsvg7d+8E4yorRrDMyOJ9/yxFg37+Gke/Dy2
WRi4SVGsfJ4T3MevwEreybFqFwhwcslpKP9DwDIa2klW+nJ7hXLuBJ1nBx5yXMQyLI58GnqOthw2
yFsM0yjZrqSgj75rdvzkf28o22z5wgH6qyNXgqUYSfLQRPkJxu6sp9f7NAEdBKcKgSzDaEoKzm45
R7e17CMigAu6pj1aREOJ9FH7rSZCEYlA4gTPWNwiW13BcURUMw+ZYdL4YrUX3iAB1Tcb6p4nCYTg
+OrUko1AzocOd9HFKylxHbzLeySBCPUZq+vY2qlowYagVae+Yu4f8xEyWFrs4XMtF/rZBp3SCvGY
E525fYNGeT4mPYm208devGZ9GR5+tGxC6hZNrilgJ2SEUXGNfDIDyqYdas5XVqqmSs+/rfLWucuS
PfPOikaLWsMsBvx8AW0liRJAusuKUrei9uN1a5il4cNWWyea6ERlnpD2d5ykypuhEzla8RGmDglI
Uwef0W9A1cdfn/P2bSH/URTOt89CRXj7+Gwkv2+cHplLlcEQ9DxohpT93Tgt/0VEjVCfvuO4ItTj
JRmDAqfCI+gcKISdVHLHbHSXTH3w+97BCW+bNFj6iDH4RKNhZXhG+Xb7Uu6hG9qArQi08Gh35UxP
n2c3rxvX0xzc+6J0IYJ2pMBNkWoHHGxKXpHY50NjCXmG1XQ96my4LCScqcI2wVrzwxSuTKn9nBFI
2ruH1IIuQS+01G4yifXd+VA1/gUKmSG/D3OXo/LDcn730WZhY/XeLlCxwflHxgcDIAJFbbDlRWJr
qOkh+1YMkMz06bCnIu9Fzxa/Y/vBGp7JCWqCbJgw2PBPDJEodxal9xa97X1G86vMWsrrjTXxga4n
N3fLHpRDxHPI71MVcUx9xMMsOJhrn8H/ashLpM8EFokWijSPkZRlzlwzz/Uj4khXXCckXolxXiX9
vDJMf6tWU1XW8huJ959LP/QUxGZ5UFOqABN4TF3Ew4WRaXcm4WPnvlA0oWgXLaSlH12vgtx9dCs0
uyhMue/glfOsckuNLWL4FxwKSzxlgeXUdiV52Y5NDl7ulQRALTwAf6xUJ+eOPOYloR5Eka+gLRKe
bIsgGSDfTLF6+oNz7wM0RT5wOani26afbb4DAd7meomAo2eT0i5J3owt61FTBBpn0BkIinkLykFV
NVJ0sQBOV6ptNdqeGH7POz7TaG/MiTQvmiCpIjJvfjF12MPTz0Qx9NMZ5/iI1nU4AnZ2/vg+UAo7
vDL6WrARoVGXAj5RGj9xrde7tsSuhEnHgnFDOpME8akXjiMwUpjOcOQR36AMACw+hKIx83HfV/yy
9IGr0xhTfeygVSNiQj2QKvhCeJ9O5t4NNWf5yWAb2EgnnSKdHjq5QXZx72ISXxssDrcVcaI+5/Yw
0oPqZwjuKOVI6f3Javmq57HOUkGSYsSQ8qxgOeyu6YKghpBd+QzbrJxABjMeYEyeIU0ckUWYvHhk
c7QppFN4hDtT2OBaTfYne333qcW+h25yLebNlFnyC5+zVAdxc/LM7K+5m/IGyf/hAzwwD8j9MDQ7
Rp7do3FkDQ6JXdEx6ZQTPhTh/ipnYobm9D0uWhzNZeY1os/KJ8k7wF86d43vleTedKh/nxpcMF2S
Cxx7RA68Xm/w7r1W5XPFyhlE0i6Jp6urqGfyV5X9IKLJNS9qqthmRlmLanrSV+kXgVnOoX6F2AYg
sjeQwdDkPVttPM8EWuHEkNYVjQ66ZSHIhRFFCTZSyjeNs38dpv5tmERcwKSrDk3fo3HwspepQw3j
0L1WZYIIUBaFxra4otTPDlZlCS+sTc1QivFEZoheZQK/fczFsg+HquwePw60hVu0f+VrQW6xTlDL
p1hyrL9zAwhUc8v3Y/9r5lUmIM/q/GOCvrLA8Ea7kBma+QOXbK+0qhPGZge9Ys7sVIFS5UrwaTVr
UzZq328GKMhvQvO27H8QITuV/xkoarQRFZ+TWqbgczWukO5YCoDeeZSFpHw/Ge78kb7r0dk4gzvk
OhdpigTjXIATPZCY13hkIJ2xNdfSUZ8moAbI5NMJcFAn2O2MQK+p8e7JCIiKEKcD1xt1YDFNJ9g0
wXtgIKSiDqCsfYBKfDlkpIV4PYBHCxoEslHZ2xvoYHYxGlYHNc53qu17iZJFDmqcFhd1QSTGzoj0
IH5jcTQSJtR82x4C8ao3GV7zNkKWBoLDz706sGCh8oVFwUY3hw4gcKXSARzqPLnE55y+CYWajjOx
71sDj6FbizdSdiSqo3Xdj1iQJuCNjndwsrVH0eI3K7PuJgsM2DhwWKilJz9LepgPAZtkr6zjHL+g
q/tO60PmPGgcqBf2NazvST5OJFJmFJi76V9E2JC6QATPT0NsAIP+Exl0clCjzYFrWb4dn8E8+Ffz
6hkTfogh9iBi4StQF5xc1fXF6MwgoOm12DxkZ4kr6tCMchysSoM20WwK0gIQUJDxB3316d9gsJhR
42my7gj1O1YhmYnbnZ5Acrv5vDkFo4KfNh5WSjKD6o3nxl1o0/vjuQyVUTwRuymW337ey3XIBmRO
j0KYzlAEvuV2rcSK0LvbOIhEEkxYfYwyrOTfXf4ZMzsWsidCTz7tRDh411M/+mRXZ+bxLOeVQDxC
wyp1x4balZEOz0v03FWI4PSV/ear1R2N6gXGhCwetgWhXG61WWTPtZG2mhajiAJd5oab4ijU0GMT
bhDYFqc6lPzATkWMX4EoTF56SspAF6qdl6Yzo/0yCrIwxjfCAlNK5kjU9uKzpobEcLvK/dBF/Zjs
8UkWDA3mLrjxytMKmueOvEUQ0HMG5Iacz8oVTZclO8CAUVkov7OZ4X0Q8VzZB1YCHgzfQvvd1jSa
o2OX6HsTkdmob2PU5g2H2l1uYhDkGMvGBdixjKtmvFeHCsFlrA08MJeyC2dbTsKpEX9gfLFuSVCa
TXNwkudxH0l5nDOF8X0U54MDYlVDYM6fxVsWSb1AXEqoEXRjyFiMs44UChbXlfGUWO+UJ7O+cvcU
vkEFFRNNKaj4ZIE6Km+QP1le5VDo33MvA7nxp669+gDfLymt/l9J/D3dW1uVx+UgQegv8knMCv3X
+uRe0HW3z15gztv5bceEXniylZTNh0npWdszN9Xf1l7cSvzIk6vxpiEXn1rJ4k4lIhWWfcXuij/0
0Jjmwm+bq5jU6uPgsZYHg1t7Ha7u5K3DxTpDZeS46QiMdQjTJ3UvIig+R9c5YKCHH/rULKbuDgJp
ui68BzrpitbVTUVQrtwRYCpyRGL2C4/KIC14ec1ZTkNUbJ3tIh+qrG1yU3ssLd7dnItECFJGMECj
wy6B+OxODmd7CecMPOMXUp2+NcLkCIebYiomktA/HjnSIruUIE1q3ImEeyW9Nqfk6V26CbEzg2Sm
6X01x0gqs38s1kRfxK7DiNShlmoXvbD2RzLLkF8qZO7rkd0QlIzFBd0CpNOn1fJnWMclHw/+PrOf
UR6kGoC2FGSW+/sdoPhqEtyzNb1qv+bhkegbOa+NIZU81QV14vzDJj1v6mttFacsbO10lhqC01Js
qvvIShfDihd6DJ30cQBKx8YBeHkAKHsksfcTU3yxypw49ufaKHH6LbrLHzrQJjm48D/aqYQnjQMO
5Ok/19CEcZpuXTB9kE4a7Lgq9eKwHvesbiuaDZ+p/IqyTT1qA8MRfM9zZSHIfBil0sRxFfi0aqcc
5sbpdRYrMMsA0pbDGjNgilHasOWjZcf5nq34H6J3dz7W/OpLo0Jp8mDHKqCNha9B7TM6lETG5YaX
mQovOxS9aoSqjJQeq78NzXsERNB3SGaUGy4OfBmJY3ghQydpXqmBezEXOg5OCjp+JtSriMWGGm7B
IkAd85aEVL/ynwnGuxUMFfI4T88aLGFQ8JXluJIL1MktAAW4rLjLrM/kOtDZSOkAZ1Yb1Djq4F5t
NiQHFXtV3WieXA4+KiQtasAZTxEs78uGDJOP/kT90erb0eCft7kyn+pA6NTtj0U9E3b64tAyggYc
JynVprquR80TERqliSkk9IvX1VkmFepwKdPFoj4ayWQ64lDzqNHMc32sh2SFhOdChi13M4yu+Cgl
AKExig6EXJYlg96/9ROgGsxaBhxSbrgzrAAZmJvxJG4q6GVNZyAJgNpxYoDg4JO4S3G+5By8jWhW
mfTHcTcSZAGBcRUwgRAM9MbsolkAzOYgrQAWRG3zBO8TJh43GtkXKdw/27MhHAeFtfiEq9YeF3hn
vEN3TIHoQGX+ZbMGT0hYMq6bQgy1MtojA0kwKfd8hgAeZRrHVY0X2pwDsPUgkd7yQnurjZM4jJYO
E119RP4DfpzR8F//UM5MB/ux9nk95zwpJIqe2XhRPJh2D6lyMRwSc2Qh4szwQ1+oMmxtwQKJCVm9
3e+XVb9uPam/K0deHgmNek8JtLFg1tCqYmd3Hx1HoH2CBrG9S9xvl8tYVnCe4aOgQ8YggaUU++L/
7vabqO4pg1PNiOumEbNnhjDX3fGV5A//oD7yfHanlVGFjx4t933cRu1NPNs9jORluyl8SNdhZSJq
hj5Brf9jjIqZrylnbl0WKi5fYBA7rSRDyV3jU0lzxlJ/7Z3aRVNWyNhbThxFLX9yx80Q/SFucmbu
IecGltIq7TPjik78MoxNU5gBezAGmphfqTvnmJFS19EPXk5iOC9TmnQwkaP9NeX5Smn6+T08hhrV
JpR1G634X0IT3CAQHJjIjXK6YKu1vYpUpsqeCi0dw9QAc9b/xzOIcZUG7y+gaUfXJ+IgDd44vBE2
Hy7TN5NQ4uCKfHccrpfIB6QJvqjbHWZ6qkXhuUVQtqYH5wEnDgMJ7xpXt41sraouH9Qn9ovbbFrn
Y/W2WvF6HDtF02+lzqim+gu6RTClmK8U0Rrtwh91WeJ+pniASM9ddoLknHkIeJBOZb6af66UjI7o
38okZpJUD/JBS5T13affJjTx8VGDYfDhQ3hKFonjeWD9IeA5a7rgjw9ksHJbLKa86UAtR2ZvUoqR
44QnDGzfYidkYM7vZ8sVGVIeKS4sJikuiUG6QCsE41kczMaG54wlWegoajVR8nZ/814D0lPtUJwT
AL+QAJs2wD88+87zT7X5WddnzdVhUzHUhLnmHxTo6OB4gF8afwHN3EacVl+PXPnM7ghzxyA6cAbN
urQRk00tC+P29auYkWH4CHBJHtmPWDpjnUnD4yPNxJ3RjrKNz95pm5CjoaSAhqH/k6qdyoylo2gn
ORzs1Ch2u0OZ8vhfJ1Y3IA4Z+1c0kwUqsCzzO/XGPg/jYXwC5uRUy7p8dBOVuB2LlpoFj3OfXt+x
DkkNoshkrWmDm+loxUhuM1hD4Gjg3uVP7sLvHsEEaZ6NtGzZp0xDBfQa1wB3ayFSOPFl+ZlEutsQ
p7zcGVvxcnbGdRot0hwstTWWzAI6RZKMVgWSEp8XjP5L402Io8bJlxq1FNVhafFUPHQRfOg7LEF3
Yg6jkG+bIJxJcKy2k0ssgCM/k/TY1iYv88BF6g2u4pmA6pTU2E/HFPdrbhZJYxxvNV/1hzyo3vP+
a4WxMqlJn61CWCD1Po78HSoJH5b9+8CoB656KTGOhYBK2FN5kmTw4FXdx5vvrkZZTR+BuYWB1i5J
7Pmey7x9be+9XuNx6ayCD88Z/F9E18cXXH+l7whQlIaUnkwaNYXuY3B5fejL0I+ym4hHjxgkgylU
uY2uSDKa9CrTRkv4lhXcTOyZg138x95jqq+OwWihitvwF6GlgAGIn0oNt9omua+5+DaP8US8A+Va
pjr/uOY4S+KF77fVJXxzgzuy0/Z2xnpkx+nsce50jGfg23izQinuyYOBJbyYY68u2d8V4/rXjfM3
sO0v7Pk5E2idPdvggw07fxAt5YIGR04DTrtvTVALVIxjvCghR5WwZahiDvtrYuyyuA4dXRbj1Bda
hxLFkoesPKTGbPIE92q/0Q8zBwZP+4uIJHrwFU0Bn1LfMpCVJLRfbvct9j8F79k2D/PZcmrmwkU6
PshwU/kWEOsgqdfQfS95KQWGzK48k7GYR/be8sdFyaQFepgwpIIQAJFy/pCrLMYjmJcOBn0Yb7qo
TR57JZn0FwhXJl1Qpk5sW5ALwq/6FhrQSahfF82T2RcVcR2WYrMVP+2RfO6oUgdxIcK0SJyFd1vI
mqQwkfTzmg0AVaQ1gkWiAAJeAFSygBtB2JzFOq7AgHyp499Np/ETi3ndZEEgEGEdp32Ow1kl4gJ8
lLHmTFJ+5TyAPhvObx5pcnci6XD/ijuj5/LR9mWTZSN3fn08PT7+PYgDYRQe0Hd2LURJtVHFx+dE
Uy4AyhQ2RAMiI8BHjOt1vmJJZ2T+mycNJY7eIpC1Ix4Y7pX8xL88pwD7GPU4h196s7YR7ITSkZYB
wQphTGEP9RMZX2iIiDqQPJJPWvJCVaQOOkk0KA9W7sXk/rpk7tNhaMif1ti/jXVIMBXdZjfBUqfV
p8AgIyZYoWnZR5/+inH2UUwcM5tCDKg0kN1ERqsVaJCgwagUo8IOCFtFtqTyMM2NLSCu8oXGdM5g
QtEY09lQQNGMIp40BJGSBKDSxFDqazugO4hSlZLmHW5CU/6NOZ4Qd1oooGjbY29TG7Nm9PSYtKvX
e44k3UkOkeo2obrikdim2CYXviyKir8kV4X7N0dfNfjPu9DVCzLjuKRjnMx5Saf8nXgK0Yjt/WZU
0sTenGv+uLrnURNz38PsbYw+hr0o7W6UJAdAOjyw+560OHx0mWT+aVoKjy4urTVh83ZTApFCHA3J
qyfJYOBu4niG9w6tPBqd5RXQ6aqjpCB/Pw/9WI4pp1RnonFJGyTQQN+kOSK5uHEyI9B0SzvZUjCE
qHn+C2kbCsOxAMkfUUquKXGgV5DuPVoPz8GLGStqbCus0Ak3NrdgYwC+pKihSZRCj1CCqaTfq77H
p25BN9iOlunzWbc1TS38xwhgeC2caUPZvLIYIQ2YgJabDMeeYroOciPxEaCMK5FNxLqY1efWxvYU
7+sPYBR5ylLQZZnuASQiMOOkbxQkME4IrV+I+xjBe0wj74dZq0SjWmrgwgQrrmij9RF7zTRnwMnK
090hTqS7vnJX+6HYZiky1j13hICKv7eqKN8ztkZHMysaBGdqcbtxJH7xsOTno+EmzGY28Bgaqc5X
lYuJXC+f5EBr2knqCcy1pZ1aaRP4IdXmUrHh6o4hvSLDRSvk3ipAtoq9mlLr2Roi7SHfxnkf2kKY
RNp83jdpPeEjb8ZZhonQf0RHt0jPfL5ayXf61oXXHl8cZQzTznFPncUX76Q8hKPVTMfyJIb2/GRD
U7Ur0UDDB1tEG2g6N8vyHyhIS3ZakVxRM9ubulhzd49RfPGAwFRvJ+6P7h2qWvM3cDd/4F1Sbsz7
RF6gxJ6eMZV/9RYxRdXmX4AZHdlwkBZTyiexmS4/aQt87OA5rkWSHCUfKBcoz9CuH+91243kY31Q
HJ6pkau0uC3iin1dggWL3oCI4b94j+JTD/eDM502arEG3fE5uY8YlSQHePY/pAElm8xnN+kSGQ94
gjba8W2OpYjx8wqgUVoeb8veVszlF5nBMKGWI3LxCwGojBZE1hppUnAPKGsJMHqv4BScZjoZQt5L
4Ctxd3Nn85WijSfJ8KQU09uFHd+u+HaCOCm5W4J5mHeQQ1U9aP/H7Son2lVGNDuVbOGlB7fWmddi
b9+5LcSWi66lc0pHfJ5ifpyMDMY9KlPMcp6HZYKXiHTemjENgcGk2qiTwzpNN8SjyHOswLbCTeNw
ZIxMCLjmB6oaFuoI0IrhIe9wmdGEMEVNlW3cZnBlTSwMBR1aMgphgcMRsgYP6Bax6uiWG3ovjA1R
lLrhyOX8gDuDDXyACYXNoRNMthsDEJWMhszipURt1jLVgnV47pDsxLjhHvwANALHLPJ8mBFNN9h5
jhQm3XsRD9uouh0d9lMxRQWf3nbmQDftGXkkQKen4bmLnDPcSMN3iZbBVTYr1i7p3v4UFrf3FHBu
ZmRai79Z+WFY7ldbtEkqHEwQ73TEeTne7BuE4YVRL6VcNDxBtuSblLZhJDcZ7kyYROq+GO76CGDB
eflVjAhJJp9/Jrv5m86NeX/TphQSOtmN5qI7QH/LJ7gnM8QlvGInJDBY0w+FvNRkk6V7mmKdv/CR
tQiIgiZ1vXszGaWNPoylNisI84LNJQceyvr8vslNqz2vQGrQnT6OPPxdGucPuAwoN+VnTKykd6fe
rCdD/+JpNKj9+yUPgshwCJCxXyddOpmdMZgeOg8hyij65VMprOgLqTNbwSlFlgQPiCsUvxEMWWGM
9nn0CoQOB2qb9+0+/5BmNqisiX9xL6yf+khAP7NGgwcC/A46cQWdJFoNIytuC6TFe5qmtDTQmEAa
az3x9c9NXP/CbfDzxh0MSs7gwulbnEd1FUMbscXvLe0Eo8SHlmyerrpCNFPubnYnRgOY8HKY2D8x
gayyPVv3gQuf0PCj7QNNdOZf7Mqc1PzC09lFzrJM5tlMbgYEa7+ljxvGRpE8EsRZ0RpzhZwU+IIk
6LTwguDuxBFMGMvGoHeCsDSZxqdG49QSXrvmknzZi58o5Bbjd0Ru5vL10U5YeSgrM3mVy1MD4aWi
bI7cKKW0W7TGL1O8Ef+R9pCzp6e8KQxnLGDFPjedQfcLuKuwpdgSezTB4pv1AdsXueeV/HALCVjR
GbjjVqJjkIr06m2v6xLE9QKHZztswLby9sIWQBw7V0G/8Z/DmcJRlM3LYy7NV7wnFGxhNbS9cTRY
90YZ0OfryyKCkk8flPp2EiUaVaf4KfyL86o+q3dngJfdfE812JtIu0hjQXjdxcIiGACwdg9BeC9B
4lCwAuiJQCr5HPkipK2ZqDrGVolXz6Y+jI5s5iKhkwNZIZFPfemF+XkiDk8YJuj7IEnhI6/Phv1b
jA8038+6oY1B+6yD0etPI7cQFbXc3UtOqt5ynrjDfYQJNxKkFhnGT3kRizAKjHlzPR8uVmdcINka
Ryb8cVQC1F1Qj8/ts/QQlG+R5EaB+Ku23n2AGxCxC+FtOvKP+p0T2ZV8K6k/KGK13QQ52J4yO+aS
HcZJ/5i/ReUccoiF9tN+FE13fY8HTzqwAysTxsvdtnzgnr+72+HpjLWQHvveiHqsnFiaQaaoA6wR
8glVKpBLo6L4Q/dFEZtkSa++0ck8i6t5/+xlRXhzpht1+aytbw75cBVNQYoZSSs2ZSJCzIj3g28l
MBQ95uq0fD5qbNa//+ErcTTDfW12lQgYV/S29qMZ0v25Wd3Q13sGKKFYTa0n6wk9kmjtB/9LypAx
I41Dwst8gKSDMgRaxJEyKjXU556WDWe4qdm5osumwZ1xtTADhV0jQ3N35ODMqRzB09i8b2Vb2gs9
ZVkZ8xbhSdj8QCKet8WkIjFJhpKNOQ1H/8pKzHkJEs3bV0eeAi9pEJI8ZhyRhdO8mUfI/8v9jpah
JgrD2UHzfBT2FsH8kkyaZlhtitnUsmz/oV1OG4hGt8o/WTGV4fyX0NvFc16KaJb8dSelKYIbJmGW
nl00tLOiKQnpJbih/iKeTRmjGVGzcF2TFsxIpePjjzlrCBHjRB1ZTeewKAwoFhnWIkbkBE4Rx0P3
pW01YXzyBdhcOrnHKE3z1Yh/9KWhuI9v3nyvwKy7NHoBP+MJcuRVGE1Ysu4KRSeoLYvMqvXY2To8
wy221usB6a99RIPzOBxK/wvzDR5a+uhy1pVTGpyBEPBFJpvNT3/Me37kiSmPkGvTxiI3kB8Q/5AD
cWQHMsMYEbp8aB0GQQVjBhFO90CZrb3XWckEaDV1xuls4aTyO6qIifEV+SkAK3UJUr+eM8ZwzT4A
qd6EUjlKckhTuU8446EQKaK0lp+rSmE+188nYPJU2uOcPIbrPfAdZZwTusVEgHPYO/01Xc295wqh
ZH4yWGrjbPsKLZL2jZRmNPq6+KsexZF8ypw/VazE4QVne//ifMaVtUPZ9XywKCzQNuQdeADK3+FH
yusOVewsl3xJxaFgMGJ1+UcUiP4m7y6k7Xef1S0ixcj0eMJYHosp3ijq+uuyMD4V3oiVhIlc97Ya
PPAPPETECOpu4RQmn0Y0crfCTdBTOJiNmfQzn+nsnSYGEoVc5gksUzlPNPtJyIqItGw7C5h0k2+/
g6n42ODxWeBd0FN9L9mZPoGCDl55G3NRI53eDaQokkoeNG3tWpUn0/RKFuThxzR0yGAdSBkqpSP4
fsNqsrBZObTkubz5pxJU3l2/XQO2HPWJUmLLlg7aZGpOiAjMJyJqjllF5+ii3Ewzvk4L4RcyJUKF
qWQEq2mGSbUMWjDePVlU/qRVS33vpO2I5ATXmxsW15A4qaLQm/sqO48dtvAk9GVjyCjOjYL06ZeY
wU/em0E4AlT/jw1+6U1O4Su8XlrwEl5mv5wZQdan8rtpbekVt2lhrIh4R7bUdAfGkjuv1ZBg8Bp4
Yj2iJmzLpjg1c25QE73A+wXUoLkgWvnnCoOTFJVsCOpr7DbMt71WUlKHkyFeyPoBePvPGO5vKpZg
U0irq8F3B57gkhcVFrWKQ5BxkPA8pfF0iIFaJee1z4Xe/AcTDzWeYwUEvFbkjMXEpbSPIWXYSNcK
33awUoPUh3p06HZ36ywkBiVzEmFWhcT/Os+bm2dg+UacBD883xBlLedXow54tw9oOX2oIveZ5Jxw
TaqH7ST91a6E5oYVNyKJetPazLrolbLpP0Fg8AYqgUsY06+/PpYSIWfR4QPvMRXpTwhixst08HRd
9waie6+7kZBxwCWSc4EexRO053Hcir2qN2SjKfzj3XqU3nAePLCBhEj9XsbH3OPrVtaLLNV77UlX
UDjfTGnsvb0ZJbjpe2Ve3Y57ArGQ0GIowz/gm6Box9vV/Tt7/peTh4gBktbp34M1Z76j6DvTn7Ax
YrTvXMniWM0jaIThTHBmCeGakv6kDppEo3m6UWQd9Wp+usSRb3Xl8Gbj4luqDvmrbw13Wvln17so
wdim7Dr54zf3nOkDjt6hoTBE0aMtOVRCpWsDUqDoYFhGc6on8aLUKguMDsU+nYtGZMqrx1A8uZfV
48AFWICqz7RIxsnH5P1od+44gNt3NhLeNR8G+ywhRNF3794y2+v5+vNCnssfaVptQoaxkhuUdpcz
2iX0l1wVMis7mCv6L4EYqisUG4jN4RfWhnQ8GExx4OGl4DusUMI77mXmcOQe4bEA9IouFhdkiDO9
urB+/iO4Fg+JRkbwZLQBjVD15MDNyeqcn1wQlA4xxLLl6/kBP9H5b9EqFvMBI7aJjU07CPTrVWXv
lHsSUoM48FmqnSEqtZk/gHBQ5sVay0UjGbAxCw6enb2ZZTHfTvbdQdubD88fDRikTiX3e4uo2hh+
kTYHJV700ICsbK0ZmMdgyVYFnpZOGgcJcEzd16N0SUzvajKvhhDgolmiOWOy5hkXS7T5xKg8iKnz
jBDUumJDNgg5t8pKt12W6tqAL0uL/NnZqUf7kI7uulZvVgrb9r3C7KbneNGKE8JwXKpBE5Rnk17A
DDP+VuYeqCTdrXx34910pFFGhoFUgFOfJ70kuPebojLiNrLno+q2n4kJkbFKoy6YH27Ow+cxuc0M
FL2TuAO7jP8qguehgJNZd2jG04cJ2CKBr+KmTKe9DPX3PyNYcJaTVeEeWpaSVGhia2/h/QxrULUG
Zbq9ZDS9rWBncpdk/KCyJ8XKvjvTQGlDYugmKXPzv9BwvNl16/q/la05uN/8WMoGtHDMW0XYgQOJ
Y01AP+T6+Me3wy3my59NSF/usBwxeTilO4bTZyhB1j5u0TejNIre27xyTF+Sh+WuL3YHIIw5quPz
e67D7L9/yWNWg9ZFJv9fi4EYufFF4xTXOSnzDHQ1oJrSXC9r5mqkZJSOuwaeJSN0rNaHioSKRY/w
kc95tqsigc02o2CBDPl5nBM3cCxQobCescKkOAHfHffuB4beBI4Y1i4xb4i/Hhzsj9bkc/Zn5UtQ
hM/KxnPPnRii245Hj7VcnXx7SJwqU31UypPEIixzZiF5t2pDJkoaerqaNSLqYBeXSN+Sk0WA+obG
WKXOY/8JfjRe82rMpggyejGub2cW4uM5Bia1na0iIAfSqSBpfZxoeKOSC+gMcq7bpTdHUidf3645
jz0njNWNSzHy1J9K94kmcqf2sr2R/aHVzF8CAR+TY4D+nY1Q14dHnMj09k61CYpQwv5q+5IQwCvH
dFtv0U8G+lLUzKz5+hrS9Je6K5iF3l60w3hktKnFNNpMhrsIF3rSuepCW1rWHRqOCNTqmST00kyD
PmGwn2Q6i8eiQ3eAnner/L48UQ1hAUEyXRhTzTgsxBNTQP6+qnHBcD40uV7tWGFYGORgAyQFUocA
zqX/CFt8D9ko/xoytihEhMpsAk1bvFS71aN3ybgrfnCujW2ObSF314ZbkyN4e9twj0WSAHNTtUZf
nvlFwnkmCfEMfxf1Fgnz9iESeMDn2hBf2YR964izIt7K8H7ys1XzxIaXAx4QDBSzvxu3b48qRMni
sStR8MNWInma9OdpI3vvzz4jJpL0R5z8LhLQ5QGPqHnGz4WCb/Hexzr1fKQ6rEZFGQxNP/tSjXz5
AOF4EPa+D2/OBOq3xGZsxQniAskFARGUrubUxPXxv/628kOWgi1PPS2l3BEFpKP+R0rZ8KjHsj1f
QvTZmWzECpF+3l74VNSmWeqaxMpFV0zkHTm9hM3oOvpLAp2TTIdDdMCkOWg14ZSFb0Ai7iFa8Utm
22fTDG6eaFub99AMOvfjfDgZyWyW86vLqWFszEFMgpiASG8TiL/BWXWXbPKZonIbVXkch9FhkZYh
3hBffSnbFHRnAuNULVcYPu82ToAQdfG3I6JN0jKMiEjZOzSg0WvGwqif/vYzwk1WNx/CstXj9NBn
bahPYPWoSVMH6Qx2weRGqs94yI6wJQjW+lePfNKUpcJpSk7fBZA6qzS7VmT9/3Iuef1afGvpu0R7
RbjCkBmg2EG9Swq+l2zz/ESCB0LSXyY016TdUWWn7izmaYidHr+hTzHZlMh57SZNbCy7Q6fDEWI1
XHraOK4TswpE2NxrGBvxyzSFkpdyRCkT3z2a84nFcQRnh4aCXIrcxu466LFIu8/k+TteRivrj0XB
q5LEKVnLJ4aLw/skRol20M5Wo6kX/ygCiG/Yicy8OPBviLZ1StWh2D0PfyAg/gu8CTR81hctA28F
VijpgER0nH6482HuLq9m/OcRTB+Vv1TepmWlp+PYDAM6qh8x+s6jTaS3A2GIWfPYmgSGjVKr6Axw
+xRHzItFYgN3zBcXbB5ie9mQhAhWHtvDUJMIVYawLcCilthpeQ+YoepVIkesY2ywdK4YK93wb4sx
8azbDbE6I+Su8N0XNSOYEidjISrassI8TVSzfMMPGkDXf398S/Wu/O2L0HgVMgBLY43sS9CwNxZi
GMCczy+hmV4QOjO7aWRnUA/imG2VQq3VvdfIBdRo/29d2q/BClS11M/8FPvHy/Vwaj4voe4U8Rjz
/kWdMFmRKLix52f1P4+yn1aKEyk5tX388G6wliTrCpNTPL2LKmUzRsbG1Rt7y50oSQnOELWJx7xO
sY8M38AiaYXos9kbEW1FUAejZq0nLFVfeTKKWaxte8gz8mJ5mVdl/m/IVZFRmfV45fb+gHpL24ZW
PZvhwJ4WRnSz5Sqt+FY1iaBIAkEmOIKZX6uAnm2i3o47Ll6SZ+N+SjazoVahbUv39Le7bcv8faw0
fqCkCwTd26LkhpePb5neD3XWWZU799jKQQsEeNvwIzl0nNJEyr4Wzrv17SIbYqBJlOyGBphw8mnq
WarQG57QHqSmuu+59wVfm7PSLFIa31y+P72Nppzlg0+97ldTCPVsT4eS+jqonA9ytyHchst19EEw
/H1RCR7/n8Gn5omQIJvYWBQAeqIBea9AyMEMIk14HsvlSSHfCDCEAZLUDKZV72Hb0wKyw/unsefc
Ls+V/A3CtLOqGDeivUfG6aKkdB2wRkP5wLA4O9pXsl0YyQNtqhfFpPWM3MF2/XHpG+7vPBT4ZpH4
lnzSU6qPYCpnWY48XYlQXRxl5q7TZeM6kynQN9mti6Pac3CwnrafQJyuA1RKMxZlAkqiDtabvEDA
gfq4rX+OOCd4gHrN2VqlUhnYtFjj+CFZnDgsQ+mD0k3Bzqcgylt1rNFyQc/u5bMD/0Xmw9htzCc7
M2NaJF28XMuC2AfZoEhf/PXdMsoW/nrMzjKcUv3nU4Q9Gam/0+EaO/BtcXUyjjlQxMuH63T9ptSW
Zxqt+i2UPC6t/pXasCsWPw8PhDlWmdGyxiL4kdfnsj5c4qCqOqCkJBFA7+pORddgzO4+0R0+50su
MyobcHPzg3oqOHfPLx8AOQvf/JCpnSnz3tJEEhzM4Ky0cJri7DBAz7CfDrUZ2+QDPe4mxnjcohyt
mwuJVVZDZzCkwReF+9TPegSZLsfBgxzH1WjMGZeSnRerS8QQEaAzMAJfGIQrS7BNlJV4AamejIL7
Z4nNXYYc4WwhiBAGes/DYiuLnx56zNjfKCmpu1MDRKyxGuJGUHfSkxjt4ehWee1Q4OIA2cXAjlYZ
Znm29ZiFWcRpNHAbJX7s7GKpkIS63Ma7BLl1QFYCydjKJYBF3HOk9Kn77f9eCwqWZu7K8BWAU8EC
BuC7n1yjUg7TF/qVNUNPYfcP/luCTXEvYQdtNkNKVmTZWqlnOWC/IY9lYWUIFfosYNHWk6U6JBGg
5OUJ2uWE392hNhGpkiNmJoFwkEfT2wGsSOnOOvq/Q+TxLu1kS3E5DBMbOYJ+/feWSziuUrYUKv+2
KTU1v4oyIvr1hn/AHQhZqM5vEgxO06vMaQvvg+ody5ZsWai4J6LtRDwZ9R2eXp+DRumoqNZyBIsD
uUHmeKgJKVlxtXFRUUCqKKjtcXwc7edaMqeRdzS+d1w/vTp3USF/nEADZ2UN7Z7/P+BAQkrv40Br
U/hijc739fJj+vgqd7VmPWvOSeg+cXi38dH6c+kBMLSE01p3+7DnmRT943NB7PVmBgzyryHtqcJl
Oy7f1OY/M6sj4metaujzw4CbubhHPvsrCOeOlDjhUGv6aWNrEEPhJdhw2bOVJ1A0keFVBIY+YX7d
CuqiqxkPFLPuOu7qDkPhd3W1+JsMhp0jCHjoMUF8P6UHo+baDZFzyBRjgoh2ndj2zNR6tBPD+tJI
BWly60xzum/ROFcOPoBrbN/IaJqRgDu1OxQ2fpusMUvHZrazTDx+b9IHjw97Sj/xIgKAtHEUutjb
R7ty894G9sbEdr7HtR/fpDEMkCbrEYTlT2qcAhPV8VDb3H38gAbbAbpmr/n8wmMG8EX5ixunHRJP
DHrHfLkPdoHNUuK+wuJUFjhCshdGdVNnQw7HbtCH2rljzvjvRzOSWjk0LnZHEXUfke6GcAtkhfyZ
bqMQy3W2T1WAGBbZcZDBS/kaemq2JiEAqSOi/cgwtJgTpqjbgIeid2b+7PgxnGcm519vNsiGnuJs
UG0TPtFXLd3RLrCOjbTvR1ay5S3/9Q3s4QeztXGtxSnuMsASbF/qTlEYzlWzBAnqVIsA9J4hrXzn
X9BRC4Mcc6WvsKJzqTsHRfjykbFxmenmi5/NH+WPfF6TJSOzwhryQghC9uk2qEx+82LoOjK/ifgB
6X3tm73GeeNNCgVuJ9Hf6q0PEo2oboDdoKDevDfoIsf2xUBRcOTDd5afhJzjQk7lgx7WpfYK/Ycm
xtK9tDJkzv0a5cR3OhJS87SxrjPfnw7jeIU/GpuDFRSYJXmCjbH25D7wd9uwccl15VP0zRKnw0Jf
Lh4uRMO9XfZJFUkz+ybB32tI1NjUNMA7M0aV3FCujLGpIr8ltdO2kE2Bmx6MdVNWJwUY0rngm0kb
8+hzI1gREHMJ8XpkkVw5a2wZq80b2PmTL5N15nbDpGXTFxSkRhzTsdzF/sXrdGxPxvaiByQ6Jk6c
aKIrsRdQUgSOfyd1wKXgw1VExEWwNgzeafIqEXMbFho5L+Ba5Or2h3cb8ZGScYv70G4dbx9STKG2
vm/pB13Jf+I4DCQ917XTUlSZw0Bz+EsbamJwBtAeE5PyQHHEDLiaBbmvEt7+795ngZ98pXHfpVW5
kCGyCpxmDS/H5DZEmnwXZatPAMavI7tdBFBHGat8oDHwcYZMhFNxsvKP8K3E+Pwo0zmpReds9vFE
xBWgbhKBJAVjUcd7EydgcIrYUpVt0TmLQ4+m8PKilcRFgEad/F5NIwPoH2UKH5lzU2e2vw6CUy6P
QaZ+mC4WjPsZYZIuURLRXLrscQVw01MN9aj6miNSmG3r+fukdZmxbUKWrzV+vtkaXdNbFIvgyPNj
Xvk2EvmaQE8T/1iSUBx3lsLrtUv1J09HSBsa0VwaeCFA0rjt9yPbBdey4lS0INwNX633jqXNAsIi
KikdEeLvxpQxPBBRNHDpDLStubQI7uW4Rhom7kgvE/U5hUL82hb1IEKvrMZBLzPiL77C3G+dvANU
EZxqfy+7WOcZNOxuApWegqaaXbBVAP4FX2sKw1GIlA68yO9QYVjbmGg2YRERGIRKt529LslmhxEB
0CUefpNiKXYawzDq6Uai9+PiKZ6TevSGrZnrsdD02DPRzukkoPhY4rRRK/COUy/2rgBlkI69MBgE
k3EmF37htUVOFFt+GX2KkUidTGqCqPs2ig95m1RAfYkZnhk/P23WAgsYtOFK9z/YEF2vUEbgHc5S
oe3dhVjffnLaxg/QpfxD8WwzaQz/9OUeef/rSABGT+wYmx1Jz2H3vBnfpmoH/A+D5Y73LIFL6VSg
BT5WlnA0MQlQGvepwvxsKjCGuqPlAgmKJtPH4LtPhUz9AbiE9OblQ2CLPGcO2m6xcSwBNbcM78+9
7LxZaBY8uRIJy7bW1FAb7i8flSS7Il900q+q7DHdAKHEIN75hwCznaHfAXeve5LGXCTfTa7Yxns6
aeo69EU7YsTP2U5dTQrVkt5NTI7R9Pz6Yag7FZhA/0aSeaWea4xAr28HE5CqNTU3UgoLewtDbHeE
xHVZCxE1amBmfbxHREhMFsZPRgAmGVj0gPLxrrw62V/C3B+35zTZxKc/UL1Xq93N0juHeQRvwAJu
pqHbHhsktK6LMq6G5kDwgC5SzFzaVYykd3bqDpV/Jet75WBuo/lYnE8IR5VRjr6nybReqTcdkoiF
0VN/xf53aWG/bKzxBoteUYcC2bwHgHunGaMiDC9tjuW5nSC5iMtKcXheecx70yTV4YXun2mUGWzQ
z8pr2Fjlbq5JHCz7gNbE0VuDoGe9E5ZVlrisfDZQp7rk//SVKrz+0e9Zvn4lrdUa1cnpx8hnPrBx
8QcV1WD8osrUzxaIZdD7vLfT6AuzkD9Fu9JuI6RgwCDHX5/1+deQEVRILS5bSqlPEuIeEcRSUsME
piWpD2dmGm5BeftfFmUPhdzEwJodfdOLHYmWXMTuBrrHeKLoKqjjgS4MkP8WouFKCmnEzVqSoe0T
90Y2zT+2bi8f1zAMnZAydxcngckDM9MB2gWwQn5YEa5F+rWg4WYy5L18c0RpePZbZLUHi265PSVK
/MoD54yQpmYI4mKECIpg9FdbuA2QuT3pt+hAnASC2xiXScGttkV526x9QkIeiuKdJDLCDPQuIAzJ
Mx0DD5Q8+SFaIR5nKZlFTip83FLVbh21OGhdmE2wt4it+jINLADGefF7Sye/h3aDfutZs4fL3DZB
5Gdhb/ZyuN7unb9U/b6GxPLnuaRT53CV7cT0NsJbbxI6fxJ1tSLauAla9LY+v4egGR5vGSdDcQ1G
QSq1ndEsS/Gs7z1UiGLO+iI4jLTe22I8uHS8uazwuLiwZ0K/GebzJClpEfD+tOFR+gENe2D/gdBl
CmldYsT/0+u0EZE0hTyYD0BQFEhLAZaYNUvCsi1gNpGPA1Qi9IPbGlBSA9oFB2zfb0I455BvLEWq
rGwy7fdJhfQiKfg31/gwOBmXtZPjoaqMHioNZyQWfW8e/IY6WjKs07x63jCSfvVrNu9ApRJ4zFph
cRx9IQw4wjH/1tnBW76nzipN5CCKFYZItofcvvkO5g4okFkCPqb26/kgBbuTA+l66cjfE4qZfgvF
4HI/X1HNd514D49P2gne8B8sKfQr5Z8bf4zYGnFKHFoULraRtQ1my6nUoOU3cLtgNzy6EcJj3opB
0XJHF0hSq5i6WQHcWXQD0G/HvkD7rQVlIRxqKQN8G28SmSnFtxw7XRHO/zqt1uIlZEqOYcpYn8VN
mKo99fAt2nXcZhog22xQld88AKf60J/w5XhpVegJ9EYWBImvIAJaSJjr3mr6onxiuPyFyLFntmuZ
qJhRaqwfXf/rWiaqYY/CrIXrsQaAX5J9iZJZcvKlOmS1YdE6c/bbnPmvjiveb/1boKWK32MkHgzj
+USIRrtIhqDnJLsJtjysiuDV/Ez9IOW4tps3wJTxMOTXVQYyHF5jjFitCQGTM0Z9xlj+KwS7awUR
XN92JQGd6JDIA4s7HPZ2z0e4DKIuby6NJrY0ue9Qvm8X50lc1UusNrv0PoJ6854NgFqiiRQRMb+x
jmNohDOOrPdCcGuCs5pnxrC129oC0csYc7F6dCFNO0DHqWxgRc2sgAz4Yq/NVck2gDw9972mdv5B
5lF5Gy9ayaQLf2+YDW/vwt9LBh+jq+5smyd8Udtw4jEO42JFtAPeoA5gaxN9GVPpW1mhVzHjcAip
C0Q4TOe1eEbjqrJGV18QSdApUW2CKhMk5KRmm+QRvWV69SWso5C1LN9AkRfob8UG5tGqC1Ov58Yl
SWlk0FJNIN7+t0E8t0FWHxn7XvjlRbPbxlJ0KE2R1xBDV3DPgFCxSX1VqqEXMlq6pD5n2pBVkA18
mluRGzUtghSuClk2Vh+HJLdkscHEB6WbQU61m8xg90TqgaqDf7VzhJV/PMEkoqsffQl/sQukpMcP
BulrBrp6WsYWqXuouCCyHt0E1fN8YgEAnEncUE9oeedJtW/dnvE0qieqfnT17IgUoqzUB66QHLGk
zaj6BcszfhFkRdo+8A78k6QVB4xifeR3cayKcBUHdKve/z6Ay62FTQf2UZacFTgZjlBjjkkx+K3Y
NV7k9dMPQA0ppt+Fo7wz3dK/BJ/wCPyXE2j4N8X7HDLnaZ9CwmOn2TrOLn+85NbGaZI/tqhRy926
iY9VyrHLi1ljRsaDiFGF1fETj8Cy29jCxLZguh4wp9aJQLlrId2Luyyj1Mp/N0PUfQM4U9oKj477
1mHWwSQ1PU8x0nX6CxmI+OcPpxP0yJDSlOtc/fxmbtJJpnKiqQLiEQyCqDGPwJ4lHNXqsq6aX4+Y
FxRR7EaTfUI3wqfiSdO1Tsa9s7FXmyHsoDu4khrRQsATEnHb/kwhI3W/SQX6AliRxl/tNY3g8CuO
EOS3WBa85tin6Gze/Vqqk7EuKS4aXAmJdvElXrGV4qhW3hZOt572dk1j7U11VNaIF7BvCrhy+E7F
Q/zjf8ITQNBTTqYCSWR7srhT3OReuVSRfWe+UMXhzQ/TK+7W8+PoQOLOOuQktj0TveJPFfvs4RJG
v2PuNfKWK0+PlTg/8DlUYlm//TPhdyOhS9dSTxaVFm/uywdMjei38WDfEP8gBcqeIl3ecqrwUmIh
NO3kN4LK6CzlfEpmXtPJnW+h4O7s2cVyNmxIS8+rtp4AwNSm009YmJXcrzJFw2B3yuvs6fotygva
kkL8EgUkjQGfqkrgScrESlXurSPvyleNGdyiSzJurYHR4oXAEmAFP6xbg8dFo2L2HmZpzfPKVKaz
v6dcyIYq27vMssrvpD7BxGjDJJ8FbqKXNblYTO5FMMYEo1pnNl0Xen3VZgmq/rLBl20o6PRZTy8V
VlikLnNoYVNBXhgLigV087NIRBIem0L4NXDjwt15ID04d5jmgd1RJSrsDRWEMjGiGkym6oyAGrUZ
glkcdy9TxDTy+HHqRolvkFNkNsjGC0ZL8HeTyqsi9uz3W3Rlma3AEAS1WQOLMglI1j84kT5h1SvF
s+rtF51NFYyQ3HoHZZjn78MVjihiK0jB5wGo3SNDBx/865ADLyFBmp4cFGyzksF6bVQaFbVKA19k
Pnfvc7eQy6AK0XaZLbfk7clBBJr1ZGoUfWMwGjrlSxsMxaUTL1NJ+Er2MSFmDNH564QNtNGok6fQ
/2JL2Bt/8lwaXVW4TtY2hz+oNgQsn4QzsBZ8fijLHf0J/Om2Mf/gkQ9J6QfS3OsHj+mbsycRRTpB
/UKzW387jtolTMi+RhrSY5gfe3aeDqEjgApQyOd3gMyvZxBb9n/X6KMB2jqbMLSFEA1c08UJIScz
j/TAHvoITNR9UuuxQQ3bAbXlo12lYasapWaRwm4PK/RyR70+r5hd3MLIOwRuKTfIBX+kANXGNqUd
Y/ytPn8z18lOD/yrFnvPpgXC4yzdm4CrD+7ZgYut114wN9Mpx0YihI6lrx5TmJ4/zXLSIsGRxbzI
r1ev2/3OujCUavthPFHFecqaMB/G8M8v8lXELeeCARKyUNutSN/vCxi8i/C29m7D8AlI2ry56Mi8
/nGBLecDkP44bnnArsH+XheJm9ixHgaxcAYWZ/NFrtiWrO9aYc/fky4I7DKEEd6oZM2fOPctscuK
+yEDIkGgioGzJwXhKvJZLClAZkug+IBXtqxMKgshaE7l788GqNbpeo8MUyruXPCaHyOAGaAsYjD4
fO+0H9rLH7T3+OPyq5QLRXhOhTd7pyOiVTickIKAFxam4a42/xm1ZvmsIYAr0+eYlzfUu7xEV5rm
qj2ErWFT0pGiX+vsXB2Q8viMbn/IcD1lW42opAMykJWL3GtG/J6Zg0N+XxCQBbeQnsiGYQUv1P2Y
f0ca8QHiE0Ecyql1KfSaXbwJC5Hi/hUAmEkYgZZnItM3eyt+EKh9VRxMB6TjAkAgyGJtiWt7ujnZ
nbv1mB6jJ9JvQJco3dFtn0jEY+a1VsdIyXkUMgVoHgir0aRj99a6yYStCR/lSTuH5FpQ4jxUyLnJ
MuHZe2127ZAghMcUF3ZE18EbzICxWFE4/H3OHkQGy5oD3P1WX+wPSwrv5cD2NxcjAMOXDUwstcPb
WEpsKPlIodU3nm/QyUsIhG4rQ6TflfvU4lnTG1K/fd1V0PJWiCJqQDxIhpYS7K6rDPccOa8irgqC
G3l+zdIDr1Rgvlw4uUM5eFZtyFIKPyYBptpMYWlggRDX59HutPZtCh7cP24XGrpP9O7tkrO5e036
ZiHJW1Q+F+W3pd/lTzyHaCXXpYSy+OKRYXsb+sLJVHZHOIefxACtI3hF8ouBdQrZxgis2IWyKXeY
A+Kmlq6Ueme0lQQqYYG66WO9qiS4mSL8fZXngqMM75Xsj3VYJ3MsV90HAHFvnLtkm/7rSekmpiwk
ltAbRjaa1n+pcfI/QOfYT75I7Itec2M0cWW4I2lrZG8jKLPvhYG/bu3KusM1ODRIvTteslGRxlq1
SGHgUhQqss1+F/Yn5RN7PupOhECMf0kyxh6hLjMl118teHf8MvlCh2gSuNTYex0URMh1geHietnP
HUr0GCQbRASD4EQffuoR4zyukIZVkJ5OAWPDqVCn1bhVsogltQSmZznsMidyHPqg27et2ubocM/2
/QKfEwpHZT01jOzVsR2jzci2Myl3pHxogoh81Oe5eyhXRzWnJ8yqElqGGCu3GEIb0NGrzU2xa/wH
0/HyHFA0cvtnUWzMdCnGhiWgT750XClfNBcwNwV4XayEVQOWj64J7iHVz86WhuKHoaTzcGOYn+KL
mL2oUVWFvT6R03OnG5IGSxfmuOe62HkV/egQUbMBK/bDx2L7R0OwuGNNnZ2xpzI2x2m9Ea3iHYW1
FM12hAZ8VrwW81pRL+eWFSa2APfaodkZG7NKmlUKebMdvEP20i9QJDAboUA2vzoTn4uloQuWJ34q
nfkIppv7B6h255akk0AyTt7OkKKINeCr/3eJBJfNr35LmzDGMgSB395W5tDfC22jVr+8lxPwOR4r
7fpmllP1io9+SRe508YHTYFPyPu0Z3vxeqgtcCAEpLWI+STDSOTXYg6gDYHeGD7FxNZf26Huqc+4
bzvaQf82OeBoqdNgbGKWn4Sk/fiyqQegtPk6jfAFNsklc3pSM23PmSs+I9UHnivO4ij1DcIk+5U7
vS6+jGUM2qwOkiO6ImahaakagtvSb99q+01xDciccjotsqbq3iHTfHfgMHsIceCl1Xfer8hGV43V
AF5trK6Jv6OuGpUfaC6BmHbbtXsPwXFQL0PgL4aacDjj5QXjDuD0rlGbHLzPRN6Be/DZU8E1RTmk
+PzOi++WhNasDYL/n7uaKK1R2FuSgqsvjg4iPwPgcbcxxn9/Byj0Cfijfyi6X1utnxnBpRvBN2p/
6Iz+Ny6UkWvhmhiYKe1blSye+m1wfKic4woaOL0XrKAXaIJJo5OPlYbnkUENiQnLa7aPWru5hJH5
y+uhKx6p2caWeE4T/GRAKH2vqlpbopTDiIiMbFRAAqZ38ERLFZ6ELhUWnEDqGX1///Z1xhZnfmvG
Pr8At9LaWghHwp6K1u4xTPI/5Yg3rDREYqltpc02SJremh+fcxQLe6Mqdojwg2ITai1ypcNVw5Jo
9ha1Pe9ogDDyLklkXn4nhNj+8ABW67VeFBy93A8ioOPncULMk9fbC/dDJrhK2Yg5heGqx4SMe4yw
sLbWdNlA5g0zQndEF7BgTnHXfaawmI3prCSYYfZnW8MPFYzCmHZMf0jPdMMrrfRVm+YiRkPZIryI
EPZIbsBbQIGGIpKpH3DLhZL61VUwlkSi3IaVbURi6bLxKkyWt0k6pZQWEbUtaDAWDFgRjvJTAFAS
k2MAbu0biVWDV9cOD2ZCqHiRnDSbPg+oYEyeHLLQorwhplz+Cy/mcq7W8Wbg2HHUhrS8bjF3hs8H
h34MxWMIW/qNs2C33EzxoqsnxpoFFNOfc9Lla3uEx8n8T7SmDQnR6BKs3EraXjIkNl8uVjmdPysw
+mwK7xOaZ3GvyZ2uaKtV5K4VJShRNHa3N9RudXrTswv8fgprsFA3ltr9++nEys92CeFN3lbBNKNt
9BViZwgLpMElYmmvxOBfMWbRKXdumYekfUL8akZB8TFRv6mkxjU4heqBwd9wiuzaUdFm9uUokJwp
9HuXhZLnaRvtmJMh8LNRa2OKyvU37AQL4xTEGPdEFB8aCCQCLTKgOGX17WFVlGVH6qxbFFWhscwE
AWrJ9Y3guyy5+cK8gIQWs4llIycAvQjRJwGyJpeiGqwmDe8BBS6P/AhTWZO/9+lMWTal5/iq3xFA
iecWP20iQqec7ayN+sY9wtCtK5rV6q3B3h2e89EorzUTUN8NUfxui0dfql+ckZlnIdw424/MwWWF
UkMJ0GgXmk3P0Jg36F4jvWCM51auhCaeiBs4fQguzZ7bPUFGzVMPSr0RC9Yhax4tOh8vbpNLWP2f
FHKNwuDgudpqaItaGF5WGp0T8p65DY5LElxn9aXgMJ43mvtRaqXRV1d6UTQBS1mZCL2QUEVeOulX
sWTKRC6nLDD/3cDXLK+9NUDG1nVjji7p34ULFcvoK6GMoakO5c8fq2v6ZaYLCfEuK+cvXg9epSX2
eixtkrdAJYE4oZh9WpfGKbriKMozk+XB6B9801n0hLntgzbJun99NvdLIsZSUAQjzc8fhYiDQ0+c
PR0vqVevp7G0iBGyXXvFXLNdNdjCIfQWYfrmpojuqwmkx8B5RcKuiEhajzdzzx5zc8Ol9tNu9JbJ
bGPpHlrw0iaOjcF5FalAnGj/G7Iclv+oM4zUPhtJWQ7+2Dm1oUbD0SZmbdX9GgklVmwkoPAfTuE3
bxlAsnFR3efmidQ12qmo6d15GPLkbOBGW/JzPsOL8KZlaIJYURkLKceSeLzaKSAtFazcWb7AQrEq
vCRmW1lvoIExofeMt5RHhTVC8egKJq3LLLXP/Fe0b5ws4DtDvcSsmBrP6PcDJUtqgNbpWSUaW71S
O9mZjun2OaLUzPqrxd4Ylo7TZH1Q1vtWaYeSJyOKJuGEQiCF2F+ccM0ALtSXEN70M9H2/m4hAMzM
hvT+okXZQEHXMoZhkoh23VCCMfifDfQxSiz+1hILRkT2sbWXEHqiJKS6rsqAPJ7iGB+mbGAWnh3j
HZEYCIl3jS32VHYaeFgAG3rKGhBj/Wx4bQCnnzRlSCbhCB7Y1sUQIEr+Z+iIohEM/cn/rHj5zuHP
1SwGXFLOI8RZZ0BtxunOYayo5Cc0NoWBk6LrQ248SmfLoYVD2O8Fe5szuX6yeoSvQ9vZhAanX+71
lw/GrNQIOdCUorPaCBSzmXL4eT6wQNLywEW+b0jKO4dumlmgzhOKGZ9XMi1BlrXaAp4BxURRt2t/
RCV16iLM3jLF6GRldI+Pnf8obv3v4f3uF27olxDxtZfKNgPxcCSyeVMl62I41zTGKM8H9/4KIQCj
WMWKxnwZYppa84l3/ihdbLzk2YJhLuRxPm7GLUDwoGD41UAZVzSlxnmJmiOQA/lZXfk7c1N3b1sf
daadg0G1Frab2jpVbWB6wfFiSckBc5VAS+MK3gWfC2xhJxQHPMYWID7Er8VPxOZOOa21g51tg93y
S15p1cMSiC/jZGfjlOU/tuJS1/sAQ4fbcovhaVD0Krc3UimNFyu6nftyqJJpONNqC7fm2XXtQ/aj
apB+h/ZYR1tKhSP/dtjYXwqqilf7pfuHt83kwVtEnGQ7FDDACRNhwabCP/7Kr2l0DK3d3C3zErWf
6gte/NxuqvhTP7eB2MnIYb2Buh0Hw++F7vt9smqgOB9FofCjeeJE3Mz2fyo/nfmx9Wk2nNYdyJNL
chBR1d/DQ5FE/VaYCkOejG+HKvNzbCKo/rlZR7GhEZ6fQTZ2NKaaXLQWcgxx0v9A+wiIAYEk6mux
3QhQgxs758s4liLv2hohiWhOWyOMl7ptS0Dc5Z2XuNIuEZ0qaffxi7eJNQsWweyUO/uwywGiGHU3
HnUuXAZPzzJxnR0AIGOGxM3bdHmzCBGS7jgiPMxZzp8U0HrLZQUUc+3x1INOmFvWIBGFOqvXHVIZ
SkKVaDNlwir8yycUUIEQiD4kBC7uAizq8wdHI2NsZrhK9EvIK4SEXIKsc7dA6T4qUxYQ0lcXhIDm
Qr1u/hON9+R6YkOc5Z6ZPwg5Qq+jEBZYif7eURNjY9p0aJfamasthT1N8VlEbZ1OkY/C6vMt3x7T
NO49zg8rPE12oWJ42+YDw3oe1zViZ9iA8JEjoGDzyWoLBWqy2KrNyAXEZuEDFmlz10Kom8Pd2tMx
E9XjbWhYvzHDh8OnE5LTJZpFo26H8yjUd1vMcOh6iqjp+Y40emXukd8q9xWLNEVMfADmH/eU8aM2
aLbmnGFCBW3rqBY5zBrNSK0/E01CUNfEm7shJoLv0Vq1fLDf7jD5o05v+Je0sgrXYwEHw4fmFv11
Qy831YdE08uAlY9+eX1Otji37TO3hujzxjNsViVd2MByMDG61zD9PaAVuw4ezs0g8R/RX+lKxRQ6
Ci4tLE6K3qW30H7E1OR+TObV2g2hxvRCR1cJ31+MaOs1Lj2vj9SyBwa1HNIAoo6+T4VdGJKroi1i
OZS1ALCm1ShxRT9vf40jWIMAdwvqQtK1S+z6s1iW2b0/IX9eG78kvprb8cjDgvoJy60qwHzIilLj
LMWDRsaBp5to/lLjVMBQ9JSgnUPOmAgJ1EGJctbfDaBRo0uLJUG/WicjY45+cJcaZr5P9qfP+bJi
DMB3ZiOedn2UZItra/c7fyNRODUhm7uWhc1n7YRgrFz4Wf65j7yYZ0wt7T4fn7aygouikT8WUGKJ
JUgt6bU2SLoM/TITLjNiYplMyGZ2wY6kRbRhIQsdsA1sHB6d/mhDs+9SiYYxpeHkQgN/hpsQpWJR
px1ZGvf9u04LNNhwTlfaBEvDcWRxP4s0ExvsxFHG0Mpg2lJFq8l0bi67MiGur51H+D8PqTNOZJJa
zfDcQc8v4e4iDg0j6vZr4m0NsQo81nb97rp4d669ZHSCtDJwr7r/R2ajqyYbT+XujgownEPSCgw/
j8MNR7egxzqFHIGLyJXz119m8vaIcxjT88TWrwjgsmL28HJSs/9N51iA9SppesWIGX/Tn/5ql+/W
XqAlZr99mie5wb0SbuMjCqDxM2l3fS1ztKFhiTsoueZkXvbPfI2fmM9DhUNzbNcWqrc0g2SXLPU7
SNTbRSOqf4/T9nyj7PD7OdJziTnXa/qtNhlyJNGa3JziTCoC3yYDc0BJnF2VRZrTYTy9u9MFHLgh
f9ZFxLjoCQ+/5AY8rlp/f3q3l6TbC1HdXOlhYl0EOkD32H5VvMjSLT3mdRSFs+gFdYUjMJDQgAQW
q5yLga6bTBAydrKxDMTAo/6L1w/K/u98evXDC5HgmEzQXOfMPjYCNKxnQX68dMqo+i7EZuBu8t6H
zOGhiXDwOU4SUoihYsttU3RJoaPci/GZEWVVnrkYkUnE3xOMd8q99SGCzimQHyyUdlvb7mIwa73k
x4oYfk1ZZt/tcmXyW3h5qdYMwwtRgVe/8o0fP/AeVAJWMSXHnYJrZ3QufpvBwhA+2PHb2V1I+YFR
2I0P7fpeuKi9Q98z0dkYIWohYoSj8H2rzgjTqTtw5sN0377cMAki3XSg95RuJyq44UGPUmnrnxf2
VQJjtq2Nhu7h05bm0xhw5pWbxGxsW6KhRlONE6R+LvgYlNPanjyBhHj5IAcMYTAsdx8xhsyO8U8v
eEPgm5NlsHYXJ+2If/fr8DuoFKeTk2Npv8n1zUnH4oweDf1rX8iVvioNrnL+FFQobE/3tpMrJ4++
XeTyHdiUOIXzD70sa+IU3PqFs8T3qeSLmVCMGg29Wlb9qFx9iaYcJegR4tGud+OSuTugBDCSuYlH
MEH0UJoiI2IErT7bg8brZazQdy/RzRanGxAmfmyyZyDw0QGKQYHempz6TXWA4LeMl6ylUh3tdF8O
Y36+NtqnuF0Ydqvze45zz90qKkOwuTm1xnEcM2aXWfqNvZkgiYdE7OYNVd096klH578k9KBoN6Iu
F4ZRtmfZt0N95vp6io/IrxQo/38fPxhYO4MW1Y+JdG4L50FwNVanfzFh7X473mtC7ZGw17HIkrXM
46MDgcLEHqqIMeWo6NJ8qFuOx+yQ4fxR3Fhr9t66opme2M9bOT+dOmPEOJyiKmRfQanxmWDq4I+M
no4FlYoxl3sOAULY3tmhtcqSJoGRuJO3xrg2okZuUpzasYkvq1Iyk86Bs6mEZIGWqV7aency1zJL
Knp8xCTI01H/lIRpNzmAoATMe2+f4Pn3j0BTbew6u24gUPeUKGF1dyPihHVRv25RyHSUHCqcD3Iv
x80yfgRB5GBCiSp8bPdDIetjT6TDTIbobT6t2JjlX1p8b2LruRQRzXQb8Tldub7R0zsHE/gew5H4
7R3EUr7lSxMhkHfkf5KieHi9Nxf1vg+npL63kEbnVPqQjScE2ZS6WDEhFQWQA1Xy3//D2G1dTctt
RS4LVHtN/3tl7fMArFkLGLAK8WKS2qOQPFbxZW11e5KF3OBHCFYsY/uUthBHnUF8tXcvvqKxmvfB
n1wH+P5HMptqCOGehjpTbz7W4DFd6eYwZKDxxRA2qnGHwTSKt6cyODsiV1B515z12T6EnhDnuD1H
+1/1QmA4STF5uAAYV8fLjZPv+vZj9yTrtQD7DwBeY/CwfufpHGqSSHC6P9yx5yNKN6rMAX0ftd4F
+Cm3BZjc5xtOKCLZdpWXgaPpZ8RJKBBBJNJp+RuWuZ/kUfYuPzpRPQ87SMJzDqZj5FOThRePYnOr
Ajdg9XJpILdLJd9ji1OZ6Yf9SgqCeoySQAcbUIbczKAE62EGxP3Q5xkeeOyQFVQDrCZZF4+s8pAI
hgm7wVctvwXBtQ68jRHkRLv3xI5O2mCINzpM4aCZX1yfERoSsdHY1Sgd0sntJQNjdm/GTQa/3tjE
vDLgqjCAWSfj6kghacvijn1f3bRZQLxlqRNJRP+qEzzp0bs5wCaFUqfv6eCBGbq6eNLZfYbSD4sw
hU0cKidaKErZ7A2+OXG5/m65hTfFtpbqg7xWV0ijO1TI2PklfmEzTeV7aVjaMxZXeYkVBr+kBznq
sWOiUVIHBM/AQDyd/HldflyzkQB6FJyHyd/fso0GHC9Je5LSGXOyPnfK2O6h9Qt/7MoWjZvsRrrL
yR66sh0FIxRyb8VwBiY7JUuZEz2TEqqorUXCEeZFBAGRNbZw6d2V66YrFIzVwauewo++YCXKS9ti
XvFXTPD6oAartQND+AUPGNcjBXJdS7AKD88q1vFFTjoAS81kf83en2iAcMMBluNWeblGs2Pe6k1x
QBPwoCyZibeQsvsSbPU1ztLbLL+veDNKMuzP/9kCTbYq4SqBnC802nCOA1+xeQ0y9+8rhCNtg9RN
MbhpXALpV+6yRynTjhfXVicLmInZjdhzhmv1t9zhhQGDKIREheGpwnw24+U+YjlFyD2mMLfUEOZ3
4fPpsi8rH9JEnJm/RlNTNlhporVE0VfRxqZui1NLYlH6w+wnAYwONTIdGUeeu46spKM7DSTZ8Pc/
768QyMzVxUYOVj7B+/x1IVu+mllUW/KnEuMP8SdrIOccd9lR0xXz6WMdWfgMOZbi39W8sKXyhMh6
p7W7bPyZXZpelectRtgGehB9I9kvdx/ZopddRYn+DAnVefpYBIxqx5YYpeJc+J3H8uhBRwHXJPXL
7WR1VSjxaEUO7Ux2rH5HeSlJPgv/jEELW9NkALvL/8295/XR21KIqPyTnC+JepRKO9GHhF+Kf9PB
Nprx7lYIWnc07AmwwTPvWj0+P2xda7f61DwnL/yiSqazkEOJu0j9lq0AgB4/P5Ndx5G2OhmIqAIR
3x0FnewPOqRjrpKmF0q7yIwZPuxMheO1Xued7Q0zxEeVSkI2/M3AzUGr+N2lbyVSAsspzvC0NMLu
Lg0ryYRX0x54sLyEwCqfmzYYTBE9sz3WGXdNiCflARtO8bvkXXZ1eJt/BJ0KWjUP4YDvbaf1sxYK
IkGbnHd6IlYABcXpoGG1UC09c90D0a2X6/RqAy/LulJxF9scrATQMMmwfat6yv/xaWi1M6Sz5Cul
jp8qE3TKsXDsxkVU+exVPuvdUQBcbk3F3H5ftgjUF2w4ff5KTeiaqhY+m1EidBBKvHFdTTcnLrCm
C4OHWllCi5t+GLDYUM3wqsUhe1NjJaY0sDTbNzTEppNbsAT0Ked/Sr+1pajRgsvcLEpiaNPlOIdr
+kxrQKzCL0Uqgf4xacLgUMPVTtE5C/PPqwAWIT/dhNH8m8OxwgJNrkflfSEf0SREq01fsdMqM+0H
qQAp0Vr7hso4ptKWl49j8biqXYzS/c/oWpPPwYig6zGPPoRBIQm48dkSGDCsr98wOodETihvLlCS
SLiJSKZknre5FJzlcsKYZo76o4QsxA8emifNY+uCqkZdglfqzwmmlfQ/VMez7hVusOn9mcHYdC3h
eZ+hoYBs5GAzPYb7HfPqBRqZoO9R/DDJj0euItdzyy6Ejk8VztTRYHAxOLRgRP+U3oOSXr+5bipK
dHghIzyFSL8sVqJT+kgdWHOuPOKulvKGvzTroxz8X1XkzhjEVGGxlrRui5QqgDr+7Qi1jYzXgb1o
5PatVLV3ONPGJBIAEdJ6qy4ci5z+1tAi3/OLmNQYBzuRolBRd/E2Hv3Pg0PL2i7iTZgpe2lxo6gF
wLCgI6JNdr8TgkcKFW9NGWxjS7Se1sxdhu9e+713fHV3jXPYWjvvU9J3kcZLB6VIvPhKa5067MBy
CdytuSpZTIMfHHd/08kgBhv/6eGfvwRsOdaoh05bPP1pOLWdij8TlLa06sVl6n8/0fO0LyiHL8Xj
bjE6SqFlkkdvux5zp6P5GwFAUNdadI3pgynoFX3GQpuXY0pGNbASfXfoUNYn2gpmGCvwxMp4mFFO
nkLZ54Lj6SaKGenmH+ZUF/YMzB8Ug/X4Bph8mprhRvywLMM9jRn0PJ18OioLBOPc8DT5+r9PHTJ8
O4tVpBuVtIocFKxbd0ypLR6Ik40oVerq/Y1zDPH4/cxqJ+oLuJ0Szy4CvYqZo6Qlgh8fj6TUrclu
V37lF4KJW4f7YX62DAi/B86cN0FH1fswsgESppwPEn5NRyGAKKGqbmFYCo+1BuI+oR1FZlBbePkf
BrLYADKe3PgtkqM4zDPPciw4su9KM4LZYjVg3yxC1V31eoJKvC3kssU4Xi+p2Vx251WVSYDZfVjI
2Q37IBbRqfNQm3O3vnTgxX2TBjXEGPkQNPMDNRLtNMpQtwTME8E0SlHcmtmtcarXKNb0/3Pl2yrb
TEOzoYGUb+GmCDh9ijofAt7cPObSLZ/Hw02PGxnNjGT0auPAo4EdycggYwjw3S/gAaUsyTAAMfpE
2akYb8G7TPFCC+8z9CYWic8OWXGWD3Ne2lzu7UR1cNrR+fTTWTSfdEcul7F1IXq3KPD6muxsX4fk
I4O8eX8PHfIfT32QnYHskgvpQk4UZ+/iq90gI4uIuvHzBpZ0pJamWo9NjBJ5ec40AnpQb6gFOCjJ
kj3UlmjsRAXZz9rMvMzRNELjPmkId6HyCk07X47npIRXDFkXFA9P9Vi7Y7uo9GhuGA8M679iD8I5
siRKjUGZFOsivwXObdTyO7boYly5p4ifsm7ZmRL32s1Gvf/jdkawsGIy5XiTThst4MCVio0RmQcm
CF9Fk6sndyhc3wu0FmM9vtjHEU8+V6V6grKmFDnDNqJtunOKx9fn6KbT/sQPLU684NsspiiC05mn
dMqfXByKkPHMfNvReXPl73CtdgQS1D5nXDhRMEhIZb7IcSmmj+Xpx102sGr5g3Lx+z+7Spld08N0
Sjv80hnsIgC0HmW5YbRSDqeAchSCAASfZB8KcJavPBnyVl5pb2wIWXHG0GJ3QR4iC7qig2hxyLuI
52XO7gduAfrepmRnBw5lhyaEnOUxCmz0b0Q3MuHAbqC5FL8MlCINOyOOF+60IJJkG0YFJLZi+Rni
hSd3dL06jdOjfQ/jik+GQFUih/kSt8Gr2pmoR0q7f2kEdbCzz3hpXsxe+zgw+5ZLBw8ZqT4CEm22
fz0y753crG5OZo0Ryw/tPltBNggFoGYG+N6mD0P29pzwLrUSGX/z//HbKsqu5nzZvloxnRJiz4vH
9zJurZEz48OGM/+SCGBm6pPWR5wYKh5XACnNEtQ5dnpBxYY+K3xFV622WKGKq8PgvvbAv0zINUTR
U9EIhARptgn0ouq/edNgxIqWyX8i2cREyC6+oJyhC2DPTpZ4eDRJiCt2Yls1saz1A02ie2pNj5Ah
KQA8e53HF4FoYn9GgZRBHNzxIBuR0ZYcbbtL+EACTUhc6C2NaWC3ba8A77Jc0lpTTCXbDF5Mvk6v
9jpdLs8xOST+c/fzCTORBymo/wS7NFbozczwG2+NezA8tKVhJ5lt3LzEySVQLRpCPzFRXAjtZqGb
PC11e5J+XC1HUNQRM53rTuculaAlBBTUdRx3HCMylRO6U8RkSiORTipiiIodFMGlDGHwGDln3mUC
wMGqECb5W7HHXJKPFYPi4vpJwWkPew9GL+5FCZaCxMp1IA+dUEaaNu85jow7Z4oy7b2nHrM2le8K
Spc9UN4/yxKl6jh05eetDbZn34pajX+AzH2jE//gkNaqdNnDLao3ZZwyhfE/jFZm8PowOgACXLPL
ZqVTfGYR9UHymnGxBKJ/5PgClQ6NLJPE5Ux9MgZxNBqOLIgruPGYugDbJnh004KH02ZB3G8cOV+q
Cv3PAeMgXd/pGmvnWUD5/GuCSe5gcKa4ZesAsNEdIot3POWWW0PivH8GRbtWYq7mugkpo8WcH9eB
QVpfrox7Kmfer08INjuA/ZU5/e3Yfwp//I4fVhbSp5YmClIfwQhFJE93lutcKaB1DoVp9dsmmCV9
BGMgMqpJT57a1/nv8g0KpWfjj+c5KZGXzMhGzusVbrp95nlkAb4p/UzH6+GPEgDxqZBCdscXtoI+
1n1VdeHrIdHoCRIT7uESZ+2onAow0AqyKpZK09KWfY5Ak1LSzN+1oitQG14eutdluCn/LekAdi8n
Hfg2p2iuPng8roVBqGzP4jIEFaqHBZSKB1+cPlDsCuBhPMSAzvy7hZQzMXSKRIC1LcZ42LTLJR/M
20zB3kyTalh3FC7v3PY1XBhaH0maB+0qW6suPfYasC+XtRiq07n6Y37yM+LPFk8NzXgFeyP71X7T
eqNmKK/aPrtgmxTPeiHyFaijdekTXpxRztGrreYtj/T26bE3gL1uy1fR17dE/aI6vzKOEZ89Z3WQ
Io8ipnmjKHTxuwGNPJ53/DN1TSh++znKR+2GKTUyk5recZE/bsHGEvT5n5j0zxDfr8B2cDcA/5kV
LJHVa/59Qf2DCggsuYOAamFA4wLpilDdqgtqOmca1XtT4OOZXvO5brsApCdMmgXvnb+RdL81KYJf
kUmPhMLP5glSiIcIH2sH53VqFAWUNa/2ig13zs5kUTFZAn2oOys6+H/k0dRXnMGdBHT/JOHUecZ9
85rCRsiVz/FoesywLzFcpe9DgrSAqAmipafjjtvi90lwo1p9Kf12FuOyevDIWQzaWB04P5+cTBMF
Ax91KBEz4TSN+SeHVffGkr+MFGp1jRsePiVgPwgGqqbm/IdLC2vvUYRZDReo8gyCVMw8dRne3dFF
o7dXfy64QwTBYFgOSiY4lfCOXRyyzTsTvIOV/ed3fZ8DqI8Bvkfa15oq3Jo8J6VwkNJp896h/MVw
1J268Y7juv6tiu/UUDO4nxY9CH+50cfLgPohmEOkApfmGZMqyT19sdLFca/AaqUeRS9Xha/fkJxv
lgKbB3MZ4Co+SAFlnTKW/ggDpOckdg4B0kmSON3gehWaV2t+hKoT756zrtBCXtxfoQq6HFhe5mlV
4YVoGoYYM+Y6qzM2oqrqsKK7o91xqB6FKeABPImldiDU9smvGWK+IPjY+6Bl1ZMuZjMNR1M+CMV7
Ws8a0zEjc3kkOlykki7j+f3x0kIKxRhB6Pfc/GSY6RgMnR7IKUMVOzNphXdrbKF7Y5HgYhRwJDWP
wzLuGx8WC6r3KQE4iO8XZABe7/wI3qQWuctv8sgm0Z9h8j+QAUjK+96udjS3JJDuctla2ldxxtOc
yQlFVOzdBbzV7JOIckdJqKHPvzgzP8oaFz8UcR+hx8FEWaL/0okGEiCqlyEV9Cto2tKjvqVFSSUZ
f0qPqRD+8a4U4bbSsOJTExmHMf7NY91qzKNrkC8BcE1mtmYTFn1hV0BTmtsmFiCPdCIcXVXRoS+b
Cuf0XNZUaVrtpf3tiNkHzUvjUOk1b4Xv+KWa77vIuMjdfq5bNiqjvKni6e6SH9EYKZW7fpd9IVh2
f5BKnqAuR4pdZnkZqHyyImrhc2+wGv7wR/1/w6CTYQ2J2I/wbPOcLqjMhSX/uZvVCOAMd+yvPpve
Wzh3oWfg+3xHG+jJweSUxWXoUVtoOWUNJnigQPsNLAhxd9FGX1M1b9ezCpN3RSUj1mDN6NTvQ2d6
Dga0gdiuDzEy0dZRaPTrf2W5bk4EABHtsnw07fWH+osr/tKlkmL60uXwr/JdKKWLLEtafLdB7hpk
DYNcTDNmeWb4ptE/0HkzmGP9rnT/uAIRA4x56qxepK7UOohtFQsrLiY2szBlD5x1Mf0TxCEna547
Zp5EN54CTzLZB8x0Tnf2uhgD1TSljQ2/PIXr4ccVryos0JzPClaL3WcIorfUHqLBJg16vJDs6KIa
Z8Mk+0sZFZ4yUvVcaI1RnyZiQ0oSTMGDLJbTsQMw8sEEnGvU7hcAHmvOw2ZZiB8/vYwXKNgzzlId
ObSh6x/7smcvXC3p7LRhgnjZgr3u0TaOaMVW3Z6Febrqecbcdzrxg32SELhIs6Gk340MYwSK6TNC
KidcRipWznrrHcoqts8L5SH89bZfdX1B5xRB4edTnnouahYQNXim4YHaM1MMfPCHX7d1XNTyYJOk
sCDVvPKuBVbsDx4Zc5FwOOgtjVN9AgApG3brk4ZnKIlJLXWJKvAZhRlzV+/P65i9mMtRvaOYzMat
U7RV2FOunubyOk0AuJAq0+puwyBBSmCYdkyLkNqnYu/mXJx8lj5X9jHO0Qf3AHRKsff97KH0XZOg
AImgPE/oGundSaeKKQquX9K1kAPaFiX07YxaURIFhx78fLfEMJAzPjvAO3IS1G0cn8RetDHrCM0t
SsHcFsbEDWYpbfRIvh6CxDN046ZtKN45A9vETuRZ2WdPJImZNrPS9tn2i3lRjqHixh5tky7MDxfI
IlcVZxEq9feiDqzP3mJkMb1Q2IIAzemK6qP9HGMTezn3F+3nq1VI7kdPgQTtTW9y1iJtlRbEJFHA
ss9cIJyin+EHqd6rY5PAHL1y9jpc8y6Q0ea6SgM7xbtwDyUoJGLNa0Sp+QUDg1/fxLj2fZQjZ0Yg
MPrlbkumIjwwVsU9Q96Z3WdLsGy8wfYIaAd+zzjswR5Z8zXfPASnVrZFZVsUV/Jq9kCYn2vN+Dg1
r6sAFqSbbOuKglv26eBH0vfukzMgJqmXfdFFBb8rhTUkSlZxzPsCO2WR++7pr5vy6vPlJ/87CyJj
QEbTDvLUqT1KRRweLdwEq+/iWvLv25EZB/gTrPQv84bS8PZ/HIRcTtKr6Cafvq+pWa4YMAHt9xaM
f1C9CKxslFPKLLNOAyDbmd5ht0mNPXPKwIkUI4vEkF1x0n4KtYt8vScg8KebUtMW/6qcZWzTvSrO
ZuD+78IqddJCFggy5Pc0jO1RjITHwqboddour7JpFj7INHoVFhySs+shX6vzCA85vbaX5utVEBIq
wf0TXDGTFfJ2lb4NeD9ij4GA/tE+XQ3WGKGCzC7k7o1XXdOi+A5Hj/BvjZ+FKsCVlmAGleJt1X4f
s/UkajJaybO4V+UGr5iWdfHrkpEk7SFUz7tJru9MuBxyeMike/tG0ERpCf+muIHrfrCDWj2Y63vn
O8Oro20wIe6w8czghjDe3cAiLs4I8H9fRSgrgj8mXUFb5Qtw4z9aIRmCOwjEz2HAkDUyWk1+pQy2
EOGoZucIH8S7fnKiw6I9Uylw2rtwoFst+3iwCLP4QKTCQx9HUzGrIGGa+orBfkcw/tVOoywWeYDM
ucK/38+RcOCVuJXfGCYFC2q07kyjQtVW5AAkSauaHHw55sfnLsymWOBH+YMZ8Nrn13AvBxN4G0SF
f2jZ33+Tvqs+BqQ1ulBxXn0FOQPB2hIS+zUEPUdRz89ofkCo7ODlpC3amNVKjHbX25MqZGN9XLFh
oNvbv3shDQMMtaUKybSH9ovZ65VrldrWuWtxJxUreJMJVrsnJMA8IIf2WBdzo899d8vsuwVggLLo
D6/fW9NtJk9XMtnqadrUSCyZTF8u487gO8MshzrCK90qj3zdvaHwsGS+IrUDYOxZk/FYZLAvjJPH
RO3oROQLUQZAwVBbTas5Nj1ri+2qUk1BDvSxDTWxc3X1jUp99u/EVb7D0oVOe0TRrfjWFr1lQanC
dOAd6X64qgDK0HGhrQQn9AYfqnKnvV5k7E1fEypJgBQ3cRXTYixi778tq2imlFQAhBg43Lj6y93q
mb/2vt6qru+vugpf/OFudthfQokn235N1GfeCJxqnquGl6FMaTnRSgdKy7GKxZEDPc7yJkOhHq7g
pLLjt/9jIOsCSIW2DIOBfNeDXlG6Vg6sUOvWg1jyNSVfgYpPv2e4aQakk50hyBQ5wigu9SBeqGRe
ixMnVlPa5wnV6drhN8+DW9JcgEF+0ogJtLDCUXRX5+BL7y90dEC2w/OJDp8eF02UzPtsfgEIyUMD
pcFyKavQ6Szg8E6YU+vR1Aw4SbPFa+34RNz4V/KneOQgB+kgXPX1NdoOFf5otKpQ9jklCngDr97A
VubcOW+e9YxqDl1rjXadZdZO+rAytUo+eeeGBI3IEQbGLn3Sdhwgn/Xsexrz8qdKKzGkKXJv76ch
mqApMwwDMoU6vrfdB0qsLr1vtWsem5IaG/gAGRg7ydo0MIBC1oyzvNjgE7LUZholetNEk0rDeg9t
iTa1flzxvQ6DKy3//Y6U41aOuxgd3mhcRMOdpLm9Lt71ET30NhibuQ1zqHswUt3cjBF+LQeObLEj
NpVhL087u46V1bQFj2LfxsFHM2305bLz0YPUxPW0i6e0cAe+IaWC+b3kmRkMaW0iCIKI10mOOiEE
A6gq4hLV6e2JJ8s93Qkq8oPGrzlm47SHKoQSiyFmyp1SwAapwOs09Oini7ibHcuX9X2Fva3Z6oui
TUL9mtyeaCdMRZjqUxAVbnr5wT7D6a8NRu1w6mCCRfhJ54aIyEIacgEEbBArDS5IKdvDJrgk5iSZ
1oicbV10BZLfKuPHa5fjzSdo1M8rO6wOSvc/xMYRqt1y3tTCElGiC9NZE/toFHoqfghpMTehKhl/
21xbX/vl2Y+jIA9IflVIeRDZXx/Fqqz+J5UBnicO8wFn1/Z15o416r6wzSPi1UqXP9Rl97YCltMZ
BM00DpBR1C70U15rHYZ5fAhGoGlxOfczBM2sJ1go6ozSIkbiinIE7K0esDNRfiIwTRijsEfMAsiN
NIBhER6SZczgY1OTT4qzjUIG9LBA5qEqE0J4tOmeSXAQqkTLZcmHKerYRSboSDQNtfZYgyJFJ+Og
IuHlAGOJ2NxB67QtjT1uu+PGFEq8ZnVUb5bhDfN+vV9yky+i35cE7KvcL1qGhvm2jlj2WZdsbd7C
b4/NYvDdYU8vwN1E6vXr0lyRiiRebu9K+Wz7RYYkhCthpPvHW/vvYNsCM4NMxkORb2csdjCBp4Dn
lLDdTFna4Z98QHcr9HJ9HLFrAxAuJTflcTMk7yLQb54MoUiEdNPuGa3U+0cdXeTwqXXFpn4lDO/j
UuKT8C/V/tG7DDSERyWt3K4S2OF6MfEHb2//jY8auLLNjveTzp/Z3yHsGbBhJF8LZlV1V2zckJje
2Ff8IGWfC8ExQQplw6j4rUNdXk1oIWlw70p9nRWX3Y/f+5UPkK4phMErVJYa5+9kwklX34yrxtxf
LuyuUuyyfR1zNTHmG8+j+E2k1KDuccB50EG1OSWvhRPnpak31/rafRoLyF8HPEOHAPOdqkbdZzLm
I8/V1tNsKBGB5LhFEnXVd23ZeL5730EbqaDBHBBa6Gv8e5TNeEl5AMjUpdG+8rTZz+HlSjeGXssS
H5DtszFZDjCXBDg4oU63n9dTiUPrbcaa1p8jr72x0SBbzmLFD951mOzvyuqcnl7qqk4eXIjFtOLP
3Fh1Ssplg6OOQWhoHdg7n9MKSPnBI/kLHkx68HsILbjUnFLSit4MS3VBFGAK2TazXJbHsCtEkRGc
yAhtW5mZ+oUCA760I6FIuJs1jif+p69am63z2eomqjYIm75lWW7M8/ykDUmlXt2n4sOMzZrvf3rd
b9iXUcXQyDxRKGZI/DC9ziv8I5SjwCG4sO9ccrd8/xXQT/PHdgzqZUb+ljtDWeQh0HzmtEO4MdxI
FhdiFxmCt/e1KW9DvJ57JDPmlp6wv4HMf9HB0rHGcPDyXDjaqnSvSMa6LpKvZSShHtXfjrmDSUzv
h3vU0HUEnbs9tjOp1peQiwcy/nsajoWMs4S24XMNIevWN8JY6VgvbPwFlZAbM8J1WsyQFyjaXKoS
+aiadhRgQvgs0IlKsCy+glBejHg9QHpO2dq7a+uBjDHQT+Vu+VHhx2/+GGh0fs4mtoj47hhH/ULW
BRE8bUjNwH/vaMk9iuBRTa9gIugyeSosWTplyXHbR0uKr3C+vLjyU7OBcmzP+WltiRFXzsX8HhhA
hK/VirbLR4k1EqUBmfzVqGsVtr6lZDodg2X0Ix52LxfOAPrT8DvgS6Wv1Y81x91EjUhxubjPWM6U
kIzqX2mWU2TVnotpFLkEv9skxqztnVqLyIw+IG04dglEVT7FuYKyLiIJfjArPA5DTA6cX1cPPJdr
l5/SLF4qUsXP39qps2MbCI+t9zO4cYG75dJQmcgyJtCmMRYMjhnY46gHxQ1Epe3JsW5cE9KuiMSn
hb/JaizmYm5wSL84kJrQlDlsTs+gk19icq8mlvu0SkoIdMQ4BwQya/dxm5H3dROPYDkmnNx1tq/Q
+11efjxPMSbeZ9nYR0qO/TbjvpWsemLbnr80o4XAayA2yDkrUKEUg3/Z/++T4trHiZvcwpXlc8lO
x52bwRJ2fsVigAeK97uAjx3pqOd7LJGjYPCh7Q7nJFTJsFYICj7S1u4sYoXh0bJLY/Bz9fnG1bLZ
BiiXaAMk/JRp6tHl2sg/hpJzPjp7MGFPzcqWQd5ZtWW4yWrgTaczEoVO+kXCDc18H+KRgqfZvgjO
40UsNNQX+KDt5gGYOv1DZcJUjj0ROE1Aul+bVwC79mnNryRU/79C7mOjJcrzSnt2wnn4rTSZySYN
wB0IA3GAHqqtvoj0qp/hC5GW2cKjwLNcH2RPs0k+oOo4bqDjaW+zO1rmKs1e2rccuzqTf+o+/YLV
UHcPw2DFvPWr3xeMiiljeZoHu35PlJuIgE+1LJAPdJ+eZTfssV16MqD8iG3H9hWSVPobdfcKYy28
sNWcNrL8FhWNpZ/pH37AQRqRWiIbcJ1ysgxg0GsEXXnpeaLTuIula0yr69+A2WO6h1/52XUfVC8T
+YMtGFL7acZ0EfVst12MPza/tYokG0XlRbL7pev7dIQpPZ0Ydrx4T4xGlMfVKsV47I6FXL+TqbZ/
D7B+ZmZpvTxSaJMa226V27U87OceYmlH/0S4KsR+PvZJDzpH7rsfUcvpzy0GU0b+lhAongf8kv6m
1a1yoMIAcsFA8+N6REmtAwOg/wWyulcwlpr+HiAycNRZ37TkIyCQZlCvMl4j+OAY90VsjBn8qVjs
WLQyYdelzn6uujeyu5AK+IPE/zj57Ry2n4rNdDqUUgCT3Zlwc9m8v9CzTXasXSKVltgZxcW2+joD
+9F9jc1TebyPu7yzId64cv42U+xVWLG2tpUvTQ7Gm0SeyGnjc74l+VLCUIwd70mDt9yMZtopRusA
hfj9Xx4eVnGyBKPOhY1xYixvCwjhhe5YvJK/lYAl/qccIkVNBZnFMb6/1pKPLNbx0VOl+UyIfvRk
BCJJTWshqoBa4iwMlX4zauWyoytZou4A1FZw24V6o2WNKwDjQNspU9aOhyNfu2OsiYMihG6G5lIq
0mKx+fc08DGmP6gTWEmb7yHT2aR2KoFRqMQE6WpZIDYyK4zK76xJ+kcd3kphSKIH4rGDm1sPvpL6
OWfSzeMa07SifVCtn6fDmCOzbgo2AhyYWFDsz8JmCR5u7x4I1/vqgj20ySPeCvTzNLIt5tZQdn2N
9OUjewA/yQ5tCnrH5P8ZEXWcbEgADVBdWC8mTBN9i7Rb2tgquo+6QK+eYQF4oRpOzBiAzbdJwdgL
uV92KLQF7xR/WN2gf5PX9hOWmZOYBYyGbdCPDE8K5EOS/LzYreueR9gOyxiCUD0Xvb23j7Q0Pa9X
lvxAPfP9ecHBt7Is+aQLJAN0AXKUouKAfZPZn5iQvwVl01oui8T2imVkBVIJscucpmlS/B/i+LVx
wE5QZLv0wMdRoqS+zp5j5xA/4awMnwWOn7qtBjZCrGV+MXL8vkrtAoBA3BDsy1fzADXelIhIkQHL
V8zf4SAoq8xIUz0JQabdT0dfVgDMKvw8JotM15IXnCymiut65kF6lm4cBH7RsCA6RQGvWKBI5YVE
ryE9H5B9prdaqgE+ilq/0Rwb/Aeu+vWXCvOg3zSvoA+WnmodUOspk5cw+UKgiZi0gozof5zts/YW
3r/JkQ1A89962420cSR73IqWk2nkkUljvuYj7YnC/eUYKxPvpNi/hRCUZc8Hkqer5JnzDd7cBOdz
vo1JD06qpKJIRH5TTtKLKL1Bsy3uJ1dtOZ5ORdTbYxf0EBMEbuInWnWuKtrDXTGEkn9qrnmoQys+
fVX4W8crxFeZ0ycytktTLIi2A20KsvTAsKHgYCeWVwBPase4U9GRh5exU5tQhMD7Apv6ERAkoeWQ
lxPdnmZ2mMtjpB+/V4oH/uYER7AFlxatGR7LqtLC5xuwXRAO163dW/wHHFzCXEYtKKs+L7e+xb/L
c3w3fi+PmQlwfommwn6V+qmj8UjOU9Ot/D1ZDFS2ySDX+vBp7u1EeBkMJMKVaxmWkfyknKnGJgpg
m+XCi/4MrAuE/13B6J6SNHdGa6q9pZ9nNCQTpmbnbrmGsMo0F/XQyOuneI9ljamPysgJ3xNIVgHC
hlPz4NPWZ/tcEvxKP3vPihPd9fTtJca17Lphz20tbICwyVA97zbcVTg0lGYAUlERopOlXgrKwVW2
Fo7+XDHgp4Tu5aMANKbJjlh/vNCiNUhNDxXgPAVeKSBBnqbJCX64Q6HaIeZ4lvDkKYWFAYRpzmFk
VLybtTRqm730QjQf4e1nnj+hosOMmo0YRIrPwnYPpqjGZ4Kx7yFjy8zpu9dtSSqg9+GYZEl9ys4l
uNloxht5xiLWKlWWSAmCxIIkRvu8Sg6zdMMZNiefKWGVd1QIx4jYiLzKVrwmu1eagnKb11RHHGdY
uVM6pqD4LZDsg1rOrNxPUdWsYynehc4pccsyAmzrJYI20suY2JHl1+oSf4dtpl3uufTDsNZQNYH0
9m7ZvUW1+jjvs8oNGV/TZVddiRZdEvcPhckO30b9enhjYSAxIJ6q2qT/OJu0HYYn03qSGv2JnNmE
kMOQgsenOEsQirqsEQRIDnJkJEjYrVB5ljHKW3UV0q3Yia+HNGwYNkWqvWnV5kXySEGD2xCYBn1s
d6vodJkDOUuc2CR64TCbYAvivUu2zcukqf/5Qr3dNMTblozdI4z8leJtoKqhh1N3C1+ek+VFAkw5
LifiKMZBGtb9fGOAil64qIi35zoaGbeBwYkF1w8FLPfzmtOnQep5ApnQLsJO/FCl1LskEBTE/RBE
+2U5ZHYFmCcdaYh13prO6qgNrDV37cqOelyhBE9RVsVu0s7rUgCqYmktlVJmAA/VjURxH7ZMKv3B
gbRZMjZWsh2lbRq6vVmi0rv6H2K4ONZjNeAmjoj0YTb0YkgalqBUL5hOt9KZN2CRz+N55NqLHoCg
WlG4sf83RGu5yLOjvMRGiPwPIKOuW5Nb4RJJUQOEv7e5PjL1RmoVM1r7XaJCIcwLYCZ/xrRMwqJj
9m+uW7G1Y0YcOvYLBrrqjRO7wWUHtcdoZWuHPBIoHVjWW45asAUoDoh0BRPzLkLZ2Y4I93tnsky6
nDyMEnsTdpNfTGALsVX5WxrZK/kk7yuVAyU0czrQ3gHKONjSMuC+vwxk+4/eGqhYQR07CuZpGTgJ
fGd5CwjPnPM/XS/NVCSyqDfBXLQcAv2cko/H17eCDdEUi1Zum5hCOiN2n39yP3qS/mPFw7ckW0GW
Rw7KTkV0xRL6c+a2/fj8sEUkLG2+5mydPNAfmIhMyMI4xoGrWKq+jWpy4Fsii1fA41dfC3pGse43
0jQLRz7GWHBruk3748C6fuFIth7WqOfBxZisXIIiOLxjbq0bXRoL3GjAQMIIStxM9xDnXyB/9Kwh
MHUAgyhYG5zigXIFA+oWfeD5ajH1tvbpixsPImaNJTLfHRBLJhA3KayeXl/twHZZUbWhXsqVZG6d
l39AT9vZzJrJZCJfUKoxL9aSoL9Xi1tj2x+yyFvNzoXzDGJF/GaK/4oWXQrpVmlmgYxfQUKaRxrP
r4ejf32rTAtM6eeJBxjHgyR1NmOrrQASlP4H/p46XmjoRC9p186ntsMjYREt99r/bYDg2mwy5Bnn
TgTwY6t+C3SKwNKg33WJquhKP89Eb8XTyDo6YXr+zNnp2x3pZtHRxuFhEPkBSli4ExgGLduCXoL/
2jWbNK/kJj9wJCg9/Yk4093m6EfhMLg8xWnoOl9N3XUwM0UxsE/Cp9QZcLWxn+xy7BfZDrSveRRV
cNJE+LqIpUiitsONPByoXOW44828AkAJTELXhVWfcrHT/qH9JESdVvzbSSKmRVMBCi/Sev/8EONg
MN/PUqlwdiZYX96jz6BGQySaJY0Ob1zhhop/5GasGWe4UCZpBL4aTjvu+C4ST93YhhuprIPKEffj
2ieHllQzWGewF4B6C4CAGPhlF2gerUjddpRQqT13fikpOJOv8zzWO+Tq9qvqdcbtwaGwuDsiUvlO
cjB+s7EvtIJPOkiwMqmF58IkFZOdsEg0nUHWP9lCJ8FDznxfr3LefDy1cYBtxQaLEAdqhg5NGOU4
8bl4YUx+EFWlf2r1HWokTGsATvam9apmK5LjXtzJfbFtUfqqcNycvP8o0PSpTa8WiKU3lx6EDJbW
FlEwP/OhLaZBqjEWWNy7+/jBQYDt1CM/5WEeXwovpo0riy+zlSd5SjCu44csBdk0NhMtvzrEZdC0
0b0EdLvvSb0/9NQ7P5ocndcHrv7KB4/X2uE+yuVdFErSrzUC1dVV/f+RS/AhtUj/MWOe5fvQC4eo
D5I7qwnfUyV16h51W260FtFR24IVeUnjvtt+sd7HTwFH5APY8O/oAwcng0RvXf0XJrFuUCVwgJvY
9jd4X4OugK8/nH/6UpNaK96VHYGP5+AnNma/YDC8ujmJTNtp7Fg5E/NzpcPdYd0xbJfMQsEXpx5d
IZP3fzX61l1PilIa5ui9vtJkyr6bqwpXt29WNqEAoJudnd71ZSGhH6BNYAr6IDjOwo/Q12AQov1t
diQOsnyT1fdvAWfRbISn4sL1X8HOCSfClvx+LdzpZCweuDzkUIw0rOQSFp8XCQPmmEHJapd0ehb8
rIYwDVV7XRWGA/89vs6NFtWK4VJkxO1v+urRNI8OzkJEo80pgQ+icdYre+Fotnsa//6DlG5xij3X
+EOveMs3IrZNVvnHXpy/oTtK9fHpZQ5CjxQZxCdanNAe15jRWGaqekG8gEV9UCyaHmZW+2iFsrG7
ishAiFdTxgr2xQ92ttGWVLvrILv6S1CQ+zTUspPPlq2wCMOaeIy+Y9G70dZVAY91jD06pC8ns4NE
5eQY79OW4oBZvnlqBrnx0AMMIKoYO45sd1zbDBWCvAw2P0C3NrqhY32XEPRcP7TFiLv/FH6rt4nB
3hJ3H2fo6MEzxt6qUsbH+EtDRTGZrRWMP3hgHoLViHabndajCoNApO0gNH2ArxScFleYIbpAXUhp
irGhSm/gD/mhhW32WXltpVl4b6tCuBrc06aCZtmLcX807zo5PeLrZzei7FCfqpZnYC8gmgfmKlYN
BpJVvn8XHsrPAcYqKKc90YidgIL9jWBO0+SCES1c8L2RNt4V2xq86riuk1/XhO3IhuKCYkVVZYRO
SQSjMt/85VPcezHcx0/OYGElDZEMdPAQD8iLHX6JBdPAbU6tbTZ115xBAaemHOaMSh4WBnfUSL13
T7YGt3zNJoXBFLnysJB8EwU6fKrOpWdvgNMSdbWtW+rrLKIg3eD5GAO23qzgND2zBnH3EqcV0xxQ
vUYYTAu8bgnJJsxpl+29FezWvZLNMtxR4xpn4aLCCDN0jj7O7PGFBrF2Cq1+wa4eR9z9S4ffpfuA
YoV2oEPE17SjloXTmBNp0/DYh6rF5bEjztR4VOgPpHEFsSIazi3Oeq28UVppVqg9W6kMGZRmdQak
YNw4+YIwlRXdH1psWDg5W8vcR5L2s0Ad/sVckl6/sl8RJPm3OjA56/GYcnLBCM9D9Ems1Jo48R+8
8fOUuhN1mZ+iVGLp9HK0zUojF3uQ3jS/tx0XU5mFls9xdwJ10RXF+unbS94Hg4+ty++/ttjgEMsA
XgKXYnFe9c4i7XRmgNeXXHyAoXM2JtIm2H7lAeXIHdZACq2pRH6m6c9IIBey7opQCY+mqbJaCh1J
88RV1tmEP4q5er4LH0ufkZnEupJNNPKc8XUeeJ9ZR/1y/6+6ahFaRZFxsi9e8mmUVR1gRzobXkbj
Qb+gSPFroiba67YlReuYEPVOC3hNykArKNq07mE4LRZ3Ad36Krp3zpguZgqbQTUSieiup5Rxc29k
CyYzMEr509+obubgFumjfFugbNN9BW+KSQJqRReDMwj+ECP2b0qkGbjfq7sAX6aZQXq0jPecZ3I+
TyXEFjAADHgpTqdXJuOy6347vnXKmpwF6/kWzuhSkOqdLLKLep/nl3WPfTSv0oI4GG6N99i7Rjxh
SNuVlbsdI2H5NftwiBaW9YWsCKTw2IxL+XLQdDND6mMXd9eYs0Y8ISqZJrhgvDnRtkpKDQA8twLf
PVewU2605FElTdGmliX2Z0d0S/87wcwXEmAN7pWlyXxEV8IwIoNL0JsUk3DZGVaqxeBJBv0Cma60
pUKe30fBvfXoKkBqtK7xD6Ls/a65xAEZ3Lm2FUpi0CgRUBZKqWSPdQZ53K7JC0LwW5o0KUGOu8CC
yZGsiAmXoE78LQthQA+M/By5GYBlKEXDgVlyENv4h6DvE2XxWoYJZ/QyX9sH0Sl/YGJb5XyvOjNS
jKA/AJMWftIrI90bFcMI3hwlmHNe0nTLM8G9g3l7Jtnx4bBi2PnweCsr5XFD7zU4NVUqkMAzd3n+
zIZZd72M6NkpdcBX+cTh3OILM4VrAh4nS9BdYB2QsZH69OcLroJ+Kw2rrVXIcrftMZHVkfVEdz1N
HOGyosfRF7b3NFmN1LU5/JISbv32TioPziCkC7YpYwpsfqp7KKnUGaRug3Oh5XYm5Pgbd54imJV8
TJ3CCZ1jqVi/VAgkXAzOukLMDaStF0yb2UHb1lbi4hCIQsYt6Bx3iCywirD7b7PMJrHznBcmghE/
KCNPuENDWiH+grjSopL+CrDOlmWJlWvW4bJe53uE9HWHh0KQFbu9yp17wZWMRg15v5Y9JYCSNwnB
uzKSNPNQk+bXE0SdrZrOMONBKX4jIbGeUpjN9BW99D92+1MrQIBn+GRHZfknfb3TNgMKBV9LRjb3
Knu8NdoIGDEX2IPGmCNvkfcLmd3URK3TKs9cFtX7rG9OlNfs8Czj5iJfA5ng82lQB36k+0L6XPvk
/lvRbaNSqQIMo7a5t7Ar+lAyWL4+HqKzZZ1hXPZPRCKVfu/po4oYyk14A3wGteTqa0lGr9fvWs3B
pH1JIvocligkn1id8OECaK5/UN9fXuGpJoJBPnw+3vu/slfrP4ufsYZsKxVAwWPBRCNusZRjm8JP
5S8ocJUl++aa+jW2l9gj/pgM5eeGmst76b2hLfNxckCKTgNa/mysO83N5lHJ8SapJ+tEpcwRNAM1
uGPMbyteYbBfDX6v1CJwgzBLNbibuR+7R0gSiOEMvFr05kUrEvWilmOOzTy2iPv7ZssN4ewPVohQ
yygkzArvpDBrr2iDz2jgX5E+v8C4+BR+EdXmcRk9C29xTA36p9awl3kvfSiMakEfyMPTVecElDfC
uT+/2Rhb6RfXLXXyQXOTexvPNLYgQhDTO5DwWEw3V9A8lcspQrZY7vJ1lxw0LLdRfttUT2Yw+5sS
UrmDjTTYqvc7MtE2ASowqX4lyJk2XNGTN7XPIOKQU+T4vcca4PqUjGRFAO7gJJxAFWR7inLi8aYk
1hYZRmy6jHuQhm4Zwfp8lXj0qDXMWygAHzJnif3mo8D/SlevzJWCV7aoh+MVeSb6IjPvrn3nl+vc
J66TKUAz0UrAwYaU67RjcxR7IWs5hatXapQJkkTGc6xtep4xyQ1z6Lg8QfnXXfO007nIJHdzoUoj
zw+BWI4cbK4lmAUdcLbnBx2+BXI3kvrUh2J+qUGQriHVC4h34r4yBDfJtnFHaV8SI7+YvFACqPl6
+yN5+cPHUozuivCiP8hb2plKXTaNhKV/GcO0fOt2veNl+tpBTLjKTh0xb00GnlS5h8jx57Drnq4O
omgW5FBrHk+G+2T1cjmNnZDsTdNweZgRW7ch9RAe4CH0Kl6JsnKi8p0J7xwU6cnGanuismhtvFY3
kf0rb7/MqRZgd4ZAyT94HJv1x/Tx+jOiGoKxdwJP/CY0TR9emqAkbBxXY1Yj2qW70h4NfrnAj/J0
7BznNsKNph1lpvDn7TgH8r6vayHoDabZJCF45YzaIRG1Rb/xPTD0KHdfFs6MCyXyL7YHJjK5mvwy
VhuO3DEBXAUC7IXAbM/28i1z9St1oYUkxjTdOg74CaAdl/a+P+4Ve/AR1BLvx4EUQawOaEiNzlaj
hAIr5XQTOHff9ieMSxTaH7kjBSUz0APRah8SDewk6FOL2RUIFi5bjdMz92NwOLm/i8Bu4F5xUYt4
kPAbTK8GhcAJCBLjxVzcZuyVGgn/J/zFRFsGsdVemPU8KcoDGpAMbKrefhP6J2TlUcKEqGn+LAn4
dlN1cS7t8JIDeVBBUS8gI6LVBiFUPzdMQ+qXPnBLep7IEiTCw2LlR58AYRrXvFefPC9O9Wvf/Oc8
TxNEv9h6rqynYAqe5aL5zqVd8y7W3go7xNlAhy5vN7TFiHBCQyqVTXpc0QrsPsAKUxvYMXnuJ/iR
xknHI8/hpSJpiE5oTPofAVz8Pjy2TdpY638gH/Vf/IpxRx5KfVz4PRyv+EN/OPkWO8a7oer2Hz+m
wXjd4g2r/V+pmAc5Nlm9B5l2TcZKgzfhOC60sy4w98ypaToFPykR86IqNKkYfTkKCPntsCjYU5k9
joP2o9215nUKoLU6TTDPRDtQjj3TYgHXN210blVoa7AvX94fof/iULzWn3GoT29hhPiILBwJSOl0
d0/s1mrC38V6zKB24HL/dZXviANcbmZFOcMlvgGvowzu1LWzPlpfciOfa1B/K8NHeymtAv1j2ZUh
onYVNOp949Iwnqs+Nf/kAE89ifeogCOGbS7q4ETHAvPO7L1ConEVLaPQKlF23U/xp5wCCnYoSM7M
Cnwfh0OeBi8F85z18ondCQMoSvShlur+lWyg21tv0O8ePkcOfXRLdwSGUuHuQzyFV70uWvfMn/bp
zJJ9BzQP0s+1Ao+CFvKhrrxC4wBkOo8WL0VLrYmpaQo2C3jyIjKuYYYoEu7nJxbYYEADA4MGU8zK
Bn4NhCQef8jI72cdR/2FIgOlL+WVnq6MLJMsfbnKmggTOEuX+SDvzlyHCX9cZR4aSIosOObdhfSM
wePsguhOI/4vqXCAHEP0oQppXG71NCxn0ZEeWobn8yCMwefdEXIQ8R8gWJgZgqsH65X3/oKBv3F3
KKMGInpiA3sfzaK1p6867Fntd9GGM5EL+3G6TmxLs1KptNGjAvQWpzh/o+fkD061HMkPCBsWPeEi
yOuwLWbc8QDFl3kqgCxrQP17obFDwOo2F2+c0dUJSnPW3VpG63MkgSIUhhG6fYx7iPElo23L/FHW
pmGkTLw78lr5vpzb3z2k5gsZd3SmUKfD0dIM3D7jatMecCtww44oUjF+l3lk61s9AR6dMp4cawxr
I7ovHW5T7mLgdqf8qGrV+mkliUPMT6esOuaLStscz+YhO7Rzs1qticZE4w9WOhkL75qnR9hSh/Cn
ntAcoEDYKmCrTJF4+sgt2ntr12heoY/698UMWxrFRoXl0W23gp2yDge3GGxALYMMvww2GNJKt+s6
tEZXYP0bpwbcQgKXl+4vDRLVAMP0RWVs9VQSUtfganTKkdoY5AN2NlpHQXZNxcdJ3L2rKhNEP0vj
fVYX5vGi5ZbHKZ00DddUWEVxGarOOcvHUxnM19MVI8nFdoRfCrqKNiYQBXU4zlr1TUmVovcRAe2P
lOAI2hcsGItx6uBG2voG1uhz/jMq40qSGeN812mfPa3DEBrtd1e7FyKLVLPye3BiUy7AOQ2491yy
90sAIw7toodx8TBnXutteeiJgyQrXcshwEh0M5ZDqo77YvrOSrP3Vnow83+IYFWwxouCxwqFuEZf
Z2bM33VaYGy0R53OtzSy1glvyOHrVLFhHqVUOySvdEEwfhYrhVDakzREpYbC9lOc4meDHzmrPAd+
GbspnvCchUvQ1jicrw8q9E2oWsXA7rAjIY5pHPDV+WLbEUKBwlqt1Etbm8c5Opyq2NCX2VAYZYkf
Fd4qE8DNy3XNx7TMxj1B+qgQu9jpSmT8qi26Yu5gihm6QrH7WFFGQSilJ2RNNjyV5T7j1Pzw2tIR
dAsmR6fefY2PALYWdoC2q1L3iRuDqQLR0Uhl75cMG2znIs3cOxxS5yBP5ZJmOv9A0wRTFptw39/B
ETfWqkx+Zb99ee0GCsjYwupCC8OttavgsbLQq2ZfkrWt+n5iXFvtXMKkyNd/a9/iVw7Em9A2qCcS
ONdj9JzENgWN9xpjVjI5Ypjy1GhdaWlX9ZUJffqYFzXY6DeGHn0tg1asgPqYSWkw94bJQJV5xXHM
/4Y+1IDAIvyJ53J4ON6nMFVltWqcbpFNeH8u2ifxrL1IDuMtXBex0ozgIr3P8MtMIfp5eumuJbRl
LnuaaK1WuSRMskYcVXhT/VdmY8gDZlr62ueUt4QlY0nU71dCKhB3tdxVV6r5Y8wH1K+p5DEHRA8K
i2e8qb/DeKhWHO8BpftluldwnjIrdPcHaiUcPNTr2HQrU/sybcnD6DO1fU9Eq3uOEY28x+JpL35i
oLm1UI9Ad3NFy9xY4vf7wwCergxCmNY/hQgJC3iZmmoE71z5v0dBfHafmg72Sqcwfqtf9aGtjmv7
wPAVaIJFfLF2hD6GtISdRVbXvDHWCQFM8p+Gspl8NIHPpO7UaVanYWCs3bj+Sy/yjUkLJmmtO5GO
DL+Lyw07BjzRmuUh4KId+wgoy62M3aVEkb9dli8qHwzq+hGqVtemsReKLXxyIpHzrkThWwkV3dLU
8xSilDkodXQYIUfdmh89ZEU9Hx7gijFntcSeEi0lRUxE/O/qtT+f1bzgvzFdFdv1s+e0Q2BUwsgk
ShK4YU20e5D+W0uQAfY7puWRMc2Wj93i9ouDNVinCgqTC09LDz50VBkqqbwqWUvB5uY2KBPvwxA9
Xzr4kMSfcgJxsAQJrhol2vS70LtirbXACBqkGHSNd+LgqQrOtgjIpEprCS0vyuRxVUcTfG/KodBA
9N27M/RW1Ebc5kWbG+ICDwLHBkuSjr5gaToaIfgcIqjNWhfQdlc7CQvR1NEVkP9gFJh6u48sLJME
CgbJRTdZaFKmZ5hacTIB31fKWWbPK/bWp6L8TkZKA9/UCkty537ab238qIH/Fy1myTlZcvneb3ge
QRLLPpfFwQBMyJulQQqkcsCm8qBVf/TOsNQ/9p734fOTKlKQMuj2C0KlkBwjBqKUOiTMOlrDwhXB
fcbxBZGMqdHEjCofELQkZdaegXPzWs+cwQMyv6nAmvOZnl6B9N4QXTZppk2WrpgUAeNEIqCDCkrQ
dCZTGpWqj0hE7/ecBa2EOgM6pVgvoMVBCCjf5ftsa+rnCML2st91vSyMtg4fv5HOMD0Qi7wLM97y
udaK5z50I00O9TrfzzSYLJS2hup1jsnIEQB3SnVcLgoPBqTww+GxF1Ipjkw05k7J3a3MOziuVjrr
eCPci0gYGS3HdbmollFBUNhrP4ZzDHkCl8qS3F86tTUOttsXnenC+D8W5YHHIDGK5gS31YF/DoHG
WtHb8d9DugAt+szcVc0xLKUW71u8Qt+079waSnzXdVM7pd+8f1ISQ6MqViMarAA23sDCyCqu8Eiz
EIDFVRRPpEDgiYQ/6+OAB5ClwfF1Lr5BxZmfmh24TbD0I2hOgjST+xrdvEKM/feH3VkZN2R8UBIc
zJFUuLDa3joPzBAu2YmlCuXhZCAz8lNB1QpAeEIh3N0jcjqt3RgzASW/Q69GslVXV1sWMn0YImyr
HtIfAlECzsJucLsEleLgjPySn9UYMHagZrM5wx/hthjqIgD7Al1GOvcvXkhyp0ZjwzAcZgJ+wfz6
JtTjDRQUZC5MMWoUZYYU/o+U2qPuoJJ4Ao0mn8B7LQ+dWeaJqCenvPtduDpi/FdC1LhwyzrEZzOg
mtWsE+b6sIzYtO9Gytjlpcj++h/BNU0QLz4VQ3QbXBVjw6ZZ4wFD5uvmJIww/0z9WbEBqn0bovRw
fsFbIOIYHs2qu0hkJUTUoixXBF3SeI1WfI1MkWB2IDiQqtfN6ZwoTmuPNIXAlw/ZRTLgOjhxiGoZ
pLQVpb/1MDPNqYYUw4I88Z8q93pb1w6f2aX0MxUS4tjnZCMaoJwWsKeplz6fiP3r8A1A7MQMNO+i
kz4xK5U6TfxrlhoynGh47ARlYfw5zIJvj1bMe3oL5cGEfi9upWvgTuK8TsygPno3aD9iWFiwRp4U
CcmvgxvWDE8MPQibz9Zz8aKdoUeK+dNLemR0ZR5jAwRg0EC9ykVaWDNnsF4DDVArIEaWJ3YN9D/6
SGoOzOrXPD1ZLdyaYjJuL5SkARUL5sE0J9BkZcPqG0LetkqySbW+RfIhs2mxZiYpFSev620pwPwD
8QjQhaHt7I9/7IBqyz4EXlmNutv2S6zU1Jzw4Aiwu1sD75xyj6mUEabxFoPfb27GFSkWcE6FlxyZ
E/2+jcvKtbTy37q85w7ugwQqwS154GBOmzuOizsjwV/5sUQ9wc3dfe0z2/ceOqVm7kFxu1x37hGc
XhqrjntQ/tG8tFkvTNGEhjxLOQ2/dPGyR6kE07znz95QE5rSkd+Q2DngyXdN0vgcnDfwB7p1KjSz
fNQCJxQDfKphE0rSF15t0WRtPzrRkAlnRdkV7Clv4sGqI+vdZgoIvzWoc4Xyd6eLRMwajR0Vcbkf
ObSWc83mZQn6x7srUpCzif8DGKORA20khuZa5p7yCn9Q75Gwy6hxyFzlBXNWsOAsd6NCfksd0XiO
TWO6oJ18NZ/akfqtkut+e0zzowmYwhBWd1qxkYhxQZxuviCxF97cQRESCgHKfTPj7Y9hDn82uV33
sauuxQPJ5fRZdSH4rHVm/zM23c10VFvHRO7nHWWNFd1S2q0JrFpsyWG7afxK1ncO+5c/d1zFFEm+
BsxUssC5nUQltQxSmEMqVQjllCc5Zp0I5yA54mHXZAy+KIcggPuSOJ572KFDuAC71tx+qT0b13dh
z9HbyWErjeXA/lF4sHyqysbJ3d5PkjmK3XPGiNLj2d9FdglVCvimluQ90ovlPnvos52Kx+++90p+
Q0RVMK9+eLXsJP5ZptJEfHe1VFVTDiznx93+IbTym58ZH/r8h7j2qAIDGtM64M+JCUfUl87tr53J
0aOAsnZVILu2xUzYEpzC3ZZAbN3Kaz2Jb4h7HyBxgkDJkO7SWdwo67ZYHw71C9PSB1MyXN+1PBzz
7J+NjgcwnsljmnB9PLGVlKUSJfL3BMleMYsOKS530lWsEeEbdJjefGmJksx2uGC2XeK/AaamUEGi
kp/E3RTykNfa2rLscACo0HOeKhI2dmYNV0MWjRj2Bi5qr+tA9L1/n394yV0jBvVEhSB8NHllOyty
uc9ZG2E/AuksYhxsoZ8Lc5DHkCvoOXqS1TmySCnu/lQ7b/9uNA8jGnHijXRnpbFVV3uxfLuRiCp0
5WGHXX8QHxPtl8Usy95Ld7eSYoMSyndJ88naQPScPVJp/T2NpcCl2a/HT4hT3fNN76KI8sU56mtN
F52en6GW2vB800j4SArok3mjatJbw/xUO0MCkpDdK0yXKX8ZK78ndmrV0iW4M1rX+TXS+ZIF6U+I
NDxI/42Dl2Q3n+KytFD9NPiEOh8sPtFdL5SgrN6A0+2l5aQAwte9WNALWVGrpsRHIJ6kJamaqIqR
0U82jzYTcSJjV7GbQZLjqQsVwfNMAyAOefbOZJL5kOHgIBRUVGqbGb+2ZMXvL2X5NNNinWeu7Bvm
hbF9QehNbOAhuiiGi2uJAG/gVXeyvE463J9TA+B14MJkpTC6BXaMvxxA3DOMXOdiFYaD2Y9qbyg5
RmZ9sXbpki6DSE3hRUu91lD4B1rGAghtnD2QZtXl/cIifWsisXkuxCQjUHrs3A0rCdgGXXglEsz5
xl8rWV/rot0LuAd3xhO4qlsv5N5Gh6KAryeuXXpdzfwlDDtlX3OLq8lR7Os5DYD1VPzxc/O6H9Ga
IZ6OupK36zjLyODRitu94TXGDAto17Yjd4KYkIX0ieV2GUg97Gp3/zQpSY5N3qrkFNO0edvy2il+
jOEuh6vR2tl6M6EY8K7mfpi6PXJ38MG9tEt/1+djKF4jBuQ5e2uwIqR65zDIJu4OZQ2qdAb+f9ll
TG2J8suL4fu7RiXrJBPsM8UcZauCoUEEpHbthawNEnb+6tk2xoCTMOiErDYWtFwRkoKsBd4+LJDS
0dF8d4A4UCOuvjft86m/XWwgZvcy8q4A9VArKNdupOApb2BdYitBSbRv/yPI2JY12gVIb6B6a2c8
FmfYycFqj7/4z9tNPIA0f7qjrKg2vGw4xbaPu1k4NV5i1ATYj/kNIiCvSgk0Ac+uJziaEFltH1EY
4fAXRqWii3ocQJRit0/ChYnrN+Zqdd/z4MlJOPu5AtrrIZ3yZqxmImontyuuME76tBofvrdr6pPM
qWwfqh4MgqCFZMfsQP4DYzXypDwUOTtluAefq+GW7EyAAZYRCY+vBxbD93LrCONpm8fhSd+jeXWY
lO/XRVL4YIIEqPbZmbWkygL+DT4Az+xBed3sufzwNmLI07cXD6gwmCtzjrDiPom3gxh+WTo/fqkq
zATjFSecI7ZmQ7HkyhbRRJN3c9ydXzF+Gugwa7RUgtj6ivD+dj0Z0Mw6D/THeeHfkYpm+Xr/atLJ
gRNhXUokbmYoqI/2wP2ZtVGFk5OqvaW/c4xp3RhT09ut43m/gCPvksTXvLhe5fe1tbEaq3I+sCds
WLqr6lu2ZFAJesL5ni+5U1B6RkrhdD6/bOIFs053G5xMEgZU5zup5JnEJN7CGgTfGfydqOOVeZn5
3WBVfEk1y4FVliwUaAJUv5QUkSdjfBd7gVBMoQSVZVE3GiInLQfu06+tvdYkLBwkCNzkueDLFSid
Du6gOo+Rzxdq/8+6N+2wUSHXPcZ7Aoc/tgsArhrYgVGgdiZ9s5Gv9JyLLJ+z1RX9oXQ/O9BRh1ra
Zeo9pSsyQ7Caf355FLrhsvDRnzzI1dvM1oifnzxO2gjz17oPyVsn+qaa31v+vOVPKegeSRKtfosU
uhH/fu+/XTkyA1Rm9oq1yyIdYFJkBQC63zmTWCaiYlePHTI9+yvJ6UHEjfw0xoU407tUpzaC5+6G
bS4AyD/EceN8lsWdhEc9yvszimys+YkRNd9uIuHCxi0ECT8DX+F2lcjbzRgf5/Z6SYsKlLsdIJTh
98zkS8RWzzVBF6I7Kjxdn6KiPtZvznBqItpFHLgYeFwLWKVOJWYE8ickI6V/MHwHsTZGWxn+v9FG
NKnr2vGcIqH+mbbov6KqmAHcVKofcGI6tf2x4iEuqPjOHUmL3OWrNOAPL3pPI4m3SxFcOmaFEMfc
Pz9zGEckyEklW0rGhIsh+U+20YlW5lv9eqFY101ErcjYPGaC7CG8Rm1yxOlAaABfz2a1DuD+6m9h
T3Kb+OW51ktJJb6cmgPkXNFlB642hgAQDAlb+L2AliGL36D9bfcBJwMhDHV8aCQNssRkfnTRz6tq
XwFPDSip6zqHXe0AWO/Q7iQ15HFa1nZy7Z82wZOds9V5P8UEiURtAnIit1NQii1Su2eVgRFuUrmP
EGyjTDhQsSpxdR3xSDNsvfGkG99xuzcWRxpQ7nP7TkH4lkR+HE8C0SmctUBooByX+r1xWg6b3jvn
8xCTCWUXChYsTP2bkCMaZVckLkxi7J1IuItjeu2DbC3SIWeTwyqTEjk3rlNsB5X20WMONX2eP8nL
FHXlVtEP7kc/h/P8hh9Q1x8ULHAJrWZ3o3V2Xtp+IZgxtmlRbC2Wdg+YXS03mNdEqX28M3u89zv3
a97eJRhxeTuwfCTRrPRz2ymbQ1vplL5r16qTGAcyf+XCJ+OCSIJB5pfhPrJpTSFqMemvQRx67Cld
ObM2sne67V9+wIJXA4ja0FrRua7XRmKnpFRfBHWMFajq6mO7bUzP238eiV9hvdfnfjVqab03Ws1i
phiIyCtbY9PRs1mjy1Ib6M58Ch1c3uMNJhKu6wU3RGHf22IBzpXu+GnNovCdJRMStFjQC4FkJLpj
3X7JecM6x/I5js0O+e3Lxl5LmMa3TVx2eHWvd0tvQIJ3Rr+EmEq6S9KKZY5//SOoL7jqcnRGMLkp
AMuOhaJPSbl82AV0Ds55zeXbYl7q2Nj396JcvGMxVs06Vqfj6CWIxi/XO3sLPUOqlkteseMfBoBX
jWZeH8v4AFnZbivqqDLYGHtmaAWECEcMOK6pL+VOz6MTluv89aghJSmc+CCxG8QONJR6Lz0XVn8l
8cOgbdqEgWgICxa+0jn8z9lsmuSwz97UHSItRBDDdiVn71712t6/MYQKckVdZxTxVJdEn2HCnsij
G62jVvY7vgWg+TZlcHgsOxBHqfhNFZa8l+I2qcHSrAQ2ZJJrtcZtSFQKWloVJTW0BjoFab3Mz4E7
PXJ2Z5psEw1e6+/DKPOLb7bq2sseGgxkd+l1KJ4pNU3IFfKhT4dhYbZbwS+IL0dDXabPsjINKZ/1
PByE8wemDhxvOBavI63Qga4IP4cZyQuIPyzQGi+D8u/UIVpnZUmtEu62dU7ykLFIxrSeWOfzrTBi
Pvrn6vb5PMka7YkszOgpupdBmqbae8NWsML44tdBI55QqPC6nVtSWAZapuGxcydoUexRyU1YeccP
44qRFElbZkc80aJmwWU76rQlq0Q1Jk6GjG14+mep/FGJoyn92e1KXmXZ8OwRDmkTl6TQZDav35Rq
XYUwx9/LAZmo6sDt2ZTgo/aKyh7KgdtUfxh8X+L7eckaq51xqvi/M57DZxIN0/pS0yUS5Fg3tVeP
4IRdmcHYFEnVfnoXI4N229UAkw4xR5CNuZcb5k+jR4aAzEY8lPNX+51bif2SE3a59d7voH7dzW+B
Gj6Dc95czUcz3Cy4xp0NW/ppuqHx2w9M0GA/zGw4hwX7t9oSyg2OhI+lDWSQzkFF6UgOy15ETcMu
vTlJzBLW7AJeficpAoAz4xct3sEmatmGm2fpajZBMHzk5+xhy4V2Cr5/jaQ+Lqw2TMT9vOvT7nFp
aj71xmXwB+u3ZbkwuaLt64w/lTdoK67Mu5A6s5DosE9Gou6B6dBcfewY7u3wzlyo11awf33umlSS
3arnSF8AlF6PhYm3k2MYvVFRgtBHHZ8EXEmzm19tRdTrCAdOsB1NTetguE6k+sIotP9L9Cqtgrhj
M6COOH3f6M7ikSCxQwkF+7zuDsiNlBgF+m/ejH7libbjn5xZHN/9kCRYi4GujUJbEgBYH9I54hDo
JgKUV9ZlNJRPSX2KVANjVFGRghhaFyzwf5sc2Nb9uf7mGnRqfi7ITyH9hz02krHKjuphm9IAsI1W
bBVQVvbxadLngIB3nEhsz82Sg78xMWl9v/ia4WLAHFK3FVsGKIxbtX/W7sh0CQxwtlk8O/h0CjpF
i9NAdkHsFPK8K9pOhHR0LfgGrxIEPvDisSNtGTebLmDTNFo/9a5tPSsThlDzxpVibLj/fjCqvz+C
UxrA79p1O8ODm7Dwy1VBGTXiTYTb0pwdV9d+UbEsYcWR9fPjpszzwE+JdmIUiWMdiTGaG7HeFmV0
u/4Mo34zQT4P4IPVEnFHg9ptZzo/b6Cg5QXKPVaGsGGg6gHKrcpm0/5Uhf983MpadsKfcdfvQsjz
C/xU92bT8xMxOn4PmDaNUn00G2eUfmtDux9Vg2+wsJl7NvZyhfpyvSi1H64J0jGwKRO3FXq2LI70
0kOSqs53747vORZRPgDr8Ox2GOxZMFTOOCwFdkliUOHCvIuMK1KW96T8IU6S8zpbZKivwKwE7Zaz
/oe5SMEuhgDnyaA2GqXYBQVKAwTaIdk7K7MG6Kkl96Z+86DyNoV/GV3gLYHiZ56QstrMAveMD9RU
iYBXG5STPGrBamL9C+Kvj8jwwVhYcfpcBn50MsfijPeYpToVYAuKEKViFPbWNWyYC84deBzpz6Lw
GTNHmQgXqIQBndSCjEKjzijupU44F3Qui7wD5Lp6r++PDg9iQP5EP/HYziPzCGTT6EvxG3Hfn/Cr
i2aEYyxlMCUiI3HNyKoLXK4ADZP2QIrEYy+v98AGXsbaHAIIrG1zZzncaHcUUDZQQ8vruP0rfVQf
F8ArFjZWx3zRGPC1bauEEkT9GDncdhkhQa9rT/KRTkdFbujcPSk2aCDd550pHuPwHnxYys7vNeK2
kpNI+qSIs1G59z7z+QPzKdCSIsPTdQ6YTEqTuY7BHQEqaCQX38Ur4KG35Rct0z3FBNHo57zsqPYZ
HWboJ8qjyWr1KZm96XcxBmYmwZGbM0BvXAIiNzvGVJeB2SrRqdVGNihAajqPu1yOg8IhESHrqKT8
O/VD+wZgZNxzKK83lystEtql/EmLZbpC8sLxLdlponCIvGoVJdRNOofyhkw9WJfmNVVGUBTO1tD2
aY+M2nqRAwp+isS8Ase5cvGO0w5QMlFE9OrEViEIu3bXxFvNaHiaR/Toor6pXynJJZ0DpZvGokmT
lkFPVIMyMiBbK5BpRE8NSo8gppbmN4cL+cwJQyGRmn9B+f2BUByRLSLuHpimIM09/bAJzF56Vb7E
ZO/vejhgwIvUvPDnVN3ys17BUGdanv8VrEK/7RS/wdws97pG9pRFka3qP8n0IeROxsKPpdaUxiVS
zkfnTI3sHMKRwG0ggxzAG/GvyJz7uXOM1BmmwVuXzkv7IiX79ATXMIK0Dj6FIEEst1R93Snp77o6
rSMJ/vVHfOhBp0Zc3JN1ldKjXKWakUvreX+ZQs6JyjaJTcTSIBq/ZQfV8hwykPzWtQVAsyqdGk5L
mxVhwrxOaMwEwwOQ1QtdtPe6Yxb4WjAawmb4U2S+hadCtdDtFQmFG6aqIJlT7OcJy/9ZYXDdexF0
e/2+tJOzDAlTQ86N+luisJ+3/fyRK5qpyLhLKvZ3JBRIRAfd8hKV65cu66rhfERAM8Gk1vM4E1G7
z5CAqGFJfY59b7FwOyZX/8mlVxbzKz1vNssItiByzF/33J9q3uZUornFVVAl1cuiMCW7aDIBjYuR
tsh1hzMugGbb8Z6muQkufbWKzN02SbGLTZyI2Mg/MmFu3YrnnuIkTckAoir5b4CAi/TJSXthrIzu
xdlOpMSdXhx0/rnvWYS4PjhWMcGyl3hage1STYWi67UfjZfTS9PZa3mmCXM2z0g4YeyvJ+BXvDLq
KTUBJfCNonxcVAlOyniIPrIIGyScgR6WKCygE0wI/0iwcpkaZq+l0yuohgp5DaoIHEuK+QEC8r5t
6dRPHBxBswddIiNbiw8lUlkMD81xy8K7Vp8qwBtqA/RW5AlS4aP3GX4whpWkS81V0nhyMeZhWfu4
Ly5CW+sYzfmjcDXvAvGL3YITfwN23jaxX1urYK4wrkKunsQ2v9Wo6lYJW0BD/qD0LyGzTISj/U+m
f+mtWz7thhEeurCAwvxP2bXLyWLMLVDpdeHwApEKmeod0BszmEurRobVi51zNT29438wSeu3wpfr
aNSFtvJ12bflxoDfk3KpT+nbmUt22m40BTedVdnFTJbFsoz6gKRzMicDzts5QazhAclihXAFJlbb
6xF8HCzF/PKwR6CbqCIIZTAW/AuhwClpSxTjxIESLgZKxK9okZDleCRoli8Yn1upLudr43jl9inG
fFgMMxX+DLsKyVxeXbKAkvrhqJZ40m2sNYkcQVVLQc2jg4OAqkOpSbxMh5qXSVxLxGMubVs9LYg7
VXwEetlCJEoSePZSlimT8eIU9uf/7IH/8Slmy9Fb2WKL4onUBoCmhwenyiCyWHaCYZsN2v8OrAND
1aLT8wy8Xx+TwITdzZ0g3axyvyHLbHIbnDNJFrSjUORRncN6pxbITiFJNkzrR/93MTCC6jpxSP+I
ZKbCCIiNj4lHkylEJnt4pNuJ54acgeFHatbULLJtIO74rnOQw6FVJNTvuOxJbkSL5eO8b7iJLKfY
L78LSLpMQ6QtKnXM++T0cfs1J8lS6fC4VbL4ylV9RQZPa0tPTzBe9263XZ8ydX4Aps3LJwZX6IlB
VHDRUPY1hhd3DbtYjGOfoEF+M6iYcYjKCEvMXQNzQZNfpRSpLlo/pKcwhgrCp9p6kAs91Y8kGO65
x5bVNolmW3qULEsb5I9Y2A5yeU9+Q79MDFfQP6mGqBUSvDk08Mh0Bgs5FB7/BKfEVsr+/KwQZQRH
oKi2huOdf8TGuhvIFd5PnkMu2O9PYEI4k41LIXSzqw/9tbx9qpyIW/1SCxZZHavAoK1JIPwnwcUf
8FU4cn/LmIB+TP6biCU6CL6zv4/MvvDcuT4kad8ySPrwCTtYqGJI1PxuzhLBmdhARKuuV23yKyBm
sl+EXkDVOXbk1qsCjHhZibNCgienmxDlB2TOfJKDkG0anI9uqw/l0aihxvFbQgzn4LR31sNkZSb9
X+RUDFJnpQwqsp2SxiR5/7+RY4hge3Zz8S6MFfEkVeIvRtMuLCCtrXKivP5GBp4bAciuZgr5RYuA
FiOweQgmu4L++A12+a0stCpOULIWhc1yNwsGrkCYqPy7kdSUlX09CzpePk0LspqktiRobVaP8bHG
w3fzj/cVOvsTaE0dvGkDFLSf09ARmul9VqQQ/mp1oTGy/h9OmkQ7pSGRVRfp57aSZsiDAhbxNutB
8PZn4P5RAW8xCeFn1LLUWtNyh8/Wt17Iq4PFkZvyPP+4UC8Ghdn7WS3j6Nb9RUCCqx6643WFyjeF
vpWPsiF3fpgqgc1PZza5qU4wF22dB/CFCuX6JRiLV/hDdH5GZXOI57bHmgbxbIYXlCftq3435Tsv
aFf6uawtB2TfMPwBITZhlax3EVMklOYghI8DXUQlUg4+0CwVox93/HJHVRpvkzxomGSTd4LK6FJf
LmStcUoAya0BA0ET9PmiZVm5A6TNnfNelBQ8tn6IZG7uNvBRb3P+Z+pF3U0ARDjOngIm+9rcrUma
i3KbcWEPDAbMox8MXRbLR3wYzFvxaU1jACf/s7ElCG+MD8SBc+s/kI6hNkm1b7lzd07QEzev5FMD
3KTBufLecUR3o85KKWTQyh3f5m4cQT3LQE1KFDYuG42O48fp9Sw+jtVqS1ErgolQuBzKTLrj0ZDb
Un7qt8JqWX4Kfs76dfh//9TCZwz3Y9QFZKoWIfQUh72lnvRW9alColtRz0Urb+2tMlsFFrDdjQ9W
cBqlhbx6c9xD2uy5ta2rBRymN4XcwbbaIX2azuGhLKXGTnTSkrToJiAOdTv/7TDdVkDPb25taDSs
GaAxjNOTabtjHR4O07whQIL1/OcZQglIsfCCW/5tDtVLcOp4j1jDffKTMP5IkTi1ZUeLnGHLUQE+
+Is94NHaR8W2vc+1u1C9n3NigAIhRiotzUwTy/vWt94a0gXLoXqhgcx3St+ydJ+Wt+wsiifc+TGm
Ap4ntBzPU9XF7J4lPv+9l84PfJmtAd2dzkRFteRAeJmyzyieaKW6r/iTwZAXjtLzu01Yv6ad2oKa
4Ek8p0+A7ic67kbFnIFH+Jjd1EEyMnqB4jAs0r0F2MqaN2XVMHQ8zkK4fnaln1OFGUWtCKZgxcaD
wou/BbG2WNWBUC8w6cOy0mmdxkiSkg0C+30aAoVTETeK34Uhq7rvQI9U9ErRQd3lQXV7XWpRFqvC
BxOUG9AmgpL98BHWKysqU67tlEnW6REGghi30Ii1rNLZoQtqCmjjXfPdFFXoDR17RrG0vjIXfypl
pm2X0GkBTiJVO8LMK2H0RB56iUfIUjduG6th8P40H0yCVVq2ythkPwTfDAUCVfYkW8b3uUenS61G
cra5DTM76pT5BYdQW3iEEOIHAwJpgZnzNSLI5mZdSEcPFkgtqkTXbFyyTmE7xQxwM3IqSWKc7QV+
cMDNrU4DrKrEilIg9Db+nhdKVEarFYhpbE9KdEe07TXUyHffdu0593kRJYSv6ngJoZPG1uWcDkia
x1cSuh4JQHLHVznM9y5aWh9lDSjq/R4FeqGPWdGW+z5ph9DZOJ9PiGfW5Ots50qSBOUtj9OgSqy1
xzAUFjRXGHNX5vaAAsx09IoLVcBRHhCb9T+vrLpX9es5Ad1dpIepIoIUjb71cbwlvdsuhq0zdoAk
fCqU6QHVZ/sPWb93hlakBpmexqYldb7uyGVWHiJ8a+b9bgpPh1+fqOVuL/ryHzp0kdU6oU/hcPC/
ox8Zi0XnbIUfOqLxOeWgavI1PLcbR/EF8dg2d9TiHATBBB60K74Hl6lyhpRu9AchKV6PRTlebFZj
oGmX8T3N7FsZIb8WDCLXSdjRRY95YQZlvseBn4o4iF6Od7IMO1f53MJdOmk3r5sNEU+aabyiU7A9
i8abcqoWeFcbjZEAbtLA+b8KU+E8e8+4OoZkbohEhmn4nB/CSxNjQZs21nkIYsYdUBPuxCygGeh9
q2ZEzFRnv95EdgDJJkTwqy85SzjoDZzRMcpv9yBTzBOF3gXR5/BjAv5AEkG9VBhXg6gi4LHk0Jl9
CtOZ9qRTSeXwgeyHrQc5Gwgbir5ahVeSWB1Q/V6WeT9DBQB5DyeTyjG6Sxe1NJ6KqKYNpZufLPIv
ZCgYa3am0FLHuNmITrTSnq7EkeeP+ZHosBZYc3Cv0stOfcEGjlLilyNInXE5OM/KZZmjhpzH8fC9
veF3Ox70wBsSjQpZFHjra5hYWjLU+5dhtX/75oazlzfUHgFYsqQpiIXx8r+5EbPFJWVzl0Iyvble
5STcuwIw7Xm/6cjzkB2/X80pQ8JKlE0AoWxp/1e3FeUQG2LMX0lovN3Hb6bu3t6ecNFfXbeMEWYH
B0/d2Bg89oyaagyFydrM7ZAoZSZHwwEc/399pJH9QUfZNCUnL9z1IXI282c6buzGfgDt/w5BZXoH
z0lg3TpQpSEhe0BSKhGu4A9gbe1VnS7wCm2tjee5et09sTo36vhHB00QAq1hVjS3elaMpjcfR3J5
4gn12WPwFKM2tMxIsV/HtOYn2WFxfTenhqLgj3SiWM86O3nZfhXaruUuGXhqIaPNzfqmodFZsRoD
4SGXxo8vKy/A5sk5oGtBfTQihKjj0cI7C9ixfq0Eaz4zr3MheCUXp0PlA+v5jpejH0DfJ9Fs1+UO
FfTan1FFrvlSlNVGNbloCjVgeWkcFyNn35M/1qkDlDcdyuVeau7efZIT8rO9cvkCwvCb+na6+kuZ
Qg6CwC1FUf5UJm47ZtNSiFqLh+IeL0oXfrNDdeCHlQR02IerzAIGveQaARVsTV7YEuJ/Iop4JrPF
vDF/zyfkEK6BygOhrUgz5oD9KHUnv29SAbyhO2q29Jsb13Mg0f1etIDwA3ehB8rHrtTYyNIMFJI+
2+Y5RgLLWL0JAPE2hzetZL1tV8oV9RbUYkjzOW83vaxqYhwSpr/BtyDGh06Xm6IRT2hTDXLWEicZ
i6rsOVS3P5FXfc9gy5nCLvbKVMY28Zm03KOwZPjMfP17Z/yAmo7zsCmhffYw+7gEvHS4OFzpTinx
7v0O8sTs1yld0h5lPJGVKUGxibEmSgP6IkUcInwCcp/68ntiG5nf2MRftos+I9ItQvLn0GK22Pqs
+nRPz6S8hdGIu16bxgSpGhKm1kTWD2aqYt9KHzX8+LU90ACRSch3OTZyl0xm93r5qa5KjIoAOYSF
dWOrzuKuy9x3PbDBcb+650fBplsrBn79BDjyA1jM7LtiycaN7YPueOLjdp3kco0Fa414SOL5h/J2
/JRNCVapNhjG3sdUu/yZxRBiNisIDrnChWUUhrvyVi8x3ueBWCanq41o2//ib7FGZLg/tlRiQ8pZ
Dm2W7uuJJGyP8QPC71O9mjD3J8KWylXPcqhFDQRn5Yw7WlwyNKLTwnLZI9hD34zKxAsSUcc9ZQ5C
ta3/EnembCB8kFzwutDPYZoxEQmCXlMYBozgavZbVxkqOQsnFRRAjL6UDbgclmgy7iGy0ykw6KTz
TF0BbuTQ6xCMr/ZSg+TsfDX3yehWS3vk+YjcrTX/oKBuiE3H5ngmlXHjza4CHELHbT4AzYzGEjKU
NGt7RfXlH5DC3fQKJd7V+HJ5Z/Plpm1hiIf+S0G8Yhq2O7OgXBuumAx/m2fhM8yMbViWDoCSVSzP
zu4EwXSqPNTec9NV+RjQk3mmV1neL2JhinTFvikiK6+J4gZqu2Ubj1rBzxMk354uetSGq6GdOw/2
duMC/9zKQUxkaap1/wn6LQLAeBUaIasfGepSj8Cj3cHLkIrIUX7mwx4XrmDwgFVITDzfVlzJRGTt
qUFqj4D9ETS22D5nmvBs9ow9VOBkSDKnhhPaxZcW7MV4J94eDUOP64USs0/3PmCyA1fdGS3isrnC
rJgtvk28R06LeBOH5aQbrsEDODnmW0Rvr6s71CczCwFYPv9DE9SZ/mAeWSeEYESsTG5pquhYFZqC
mb3H1sPq0sMQSP130eelKUccMDuvGA2SBjKYbBMJyEpS6jK0VZwn9iVlsGsbD+KyKzkdGg2Gh+PZ
l/v/GLhIGdu/0ZKRcNOWizcWzzYAFRyT02cyrUV7PksyEBxC1AjAn0AasL5OLPyYr8g8Qy66K2Oh
m3SuvoX5DNXegWN9K/x0Gpar7zkOtOH9FedDoO6oelW1edlx+Rt+UlcROuWQqczo0fG75RTB7IZO
G/fqTOm8I3ksXyPUTUZQT0od3jnTh8pbgZvVSdz5Pbb1xqE3KckyHoTpEa0hZUtPtZTPd3HmEVXC
/iOWO1LIbvlhzmlOCsvKVCquMzSliRocLDXot/1CboumF567fW/AnCGAXQHNDTARIpa2hSH12C9z
6yHMUXZjVkf00ye2pySk3wMau9I0fgCWG3KX2k9qSlefzdeww2ySwTAFux1H6GgnWIQvjPlEQuf6
NE4y80PK8tcpHuvUtZW/pkP2OPCeskiKQpcb88uRlerqMqPdNnR7QnXL9sM1E+M0WVALTqz/w5kS
Z5vTpVP+nE8mVwbcZpLyAlapkJ4v3rcap9jR5NKPgY+DO4miItSdvZxfHiiuHj+V5aYcpR7HLMFU
goPIzZgfenYdItXog/SuUG20WbNUXgSFaKV2nNrwDWj9H5LmSrsId0zQgj+Q1G7oQyWBWRAXmRQH
bH2PRsmHVi4BoKRDrOGKH0DzeGhwuN5jSnWI6s4zHGSMyNwfReDLR1OljOP08JJbfdEFMtdayD0+
tmsVGz7z5KaZ2/YMcslix6j+Q4bTbHQK6Ev060LF/5/UKIjGLuSx2tdNjIbgWsfaryJtql1it8z+
T6c9CciCb42Z9XALW010BpEWjPGAQAgPV12GIbFgR0CXXQA0AWdJhnIU3d5f749CVF6VMjY6e7+e
93Ika5CiaQ5nbVkdSQ5j2we5vqxxefyJG8pkgEDUkxp+SFPcIXqfKpN7R0/EvWCwuk0y4UkXS5P8
T71DOYvPGSUA/oyMfYWiHothewx4vIo1+5aR7zDEvR7f0zed6w/IVdZ43qt4ExDeGUS0NY/1cZnc
uYJB+NKwAFWRwhrZmAqfkLIN9nwj5sxdjiBmByMnKN3nR1Pi00ZLSRNHaKKj0BjmZdoc6KtSo3iA
Bo//cVgUuk/sBkVcJM3rjJC84/s0phq/IJGkPMkWrqDShBI6Jx5WarcifGvJ3zdZZG9zYLUWxZ+p
ClKeBQP8U5hJQfffVjfqxt7wOGrTJwjYjoCN9hqrCuzYduTRUeDVBPqGGKly8XCANZ5MqMe62ui0
mHUOtzCD+H8DBD6c1zzahbdW5xkxNfSW6QUEPKwQ/Oo5U/LG0quxTFUCpTy2BKAMsrR8qHozNcYu
j9og3vNJDBi/fCTiS25K3VheG0c6RnR6EMp2SCPsJFRpsCxf6lxx+ZA4gUScJxpHQFboXfgCk0er
ZJ7NL2vZXTwV3lOy1sjlGh06NvFi4Pp7FQx8F19UJ22ooYVc3JsotjMTFmyl/8Nlx0JRGRooSFAk
mDlEk4KgbgsTGavuUzTSWE9XvX4lj3IfimLexlv/Nn/9C7OeqvPAC/MZ4594xJqNRRKP42Lx+Mi3
dJHo0v5ax9Y8g+tB0zrtUFQTVu7GbkA37XFsR3BqMeFpmuVRI1sHo+PuDgHA/zNnsyrjcdhAtfd7
gYqEMpdJLeRabeyPVvRJ3BnIEPD2lQR6zDhZPmt66MH56BeuqdRw4zZyNgpy0SFYazhPeNGaar5v
Q+7E3BtaItf8JQiP8PXfk4CxOlRWaRjCva1QKHZ7jcXoDh6gVQ7v9vJBJpfihtictC7Ob+iovyHE
EYRtsZI7qnM6gpU0slXLy4ivw/g8qOUsqvBinkOFD17I77p02B9Pfpc0BFd5UiHg8hOgs2muG4wL
heDexwCQgqVAmW+McfKfVlqDcf4YPEIRHtgEXTpfvkyzYsLH2BcCoIqBqtFwkMzcqhw/c0lxcGw7
5w/Ehsj9xSQhFeJnP2rkAnthFu47JtupPBIZ73PBoSkbKzKFdrBes+OIw/aY04a3Ymqj/wSkH2RJ
zVQw69U5twUonVwD+UqwTDdgubk6b2J7/wuQyU65COBvHymcaMYf8VdQZ+oonfbxavl8Bt+5mGOe
koxSoceP4g4Tdwg+38x0DLBWt5tjzRZXY7dhmn50wJ3uZfQAsCIi6Myvbv18jTBOSufEOGgH6jd+
nTUkkLeAGPbMpuvyNNXUh0kOtq2S+PjrNQXQXA5IqT4OSNo62Y7KlCqiaIn5TS5/txLgJ8qMrt7I
XMMmwv+eysYFdvUkGimSy8A7pYTf3oTSgcFQalMINRu9i/nhppxgN0gw1QwmojzEElSk8UuNjiM5
tdhe23Cfqs7MeVgBb3BC5GJoGadH4OM50B2csv0L9J5qXNYtD3mX07c+87HKuX3q1qjm49JX6ce2
yYchsZBs7HoF3o4qv7s2sr57fZRwECLjWJf0n8PFyFJG/WHOi7sxEBzTp8xXcZPQg1EJ3AoE7frc
GMeXejHFY5VHuwqPPiZU7dn8MtgpkzW42Z0lOUKnGEZQa1jrnjq5x6uEze6Fm2eFKDsYxPLZZg0H
TlhTjK7Dg8pQdNBI/EGhlDOOmUw000fABjOdrhLoXsD7jk65NA0WBwccf8ZeTsiZ582nnQjz+ngu
Rve6KH8UJMl+3xlAosh3Eo6ApvrHzglWqTG+a0ADySARB5XcK8KJk8kQ9c4rBK4D1ntFeLLMvMIK
+AMNuAveJhbP3vBJjpzorntLaMStzQQpf8K5b7Gfdll+wusZA8/1Ukqx9gyPil33XyFpa3S0WXWt
A99qxh+xnOAA+4KvS531N/eetc3rrDUViIcpiJyAp4VNJ6veTQIbXCdMe6PNMgSZSCJlNdrk1y1a
Xjj52yr+ChPcloPhYQLrf8MdxzVpPaWzc3iX3LGYoD8tRT0Xa8Ms+mDBhKBcy93k+jS3tEDDUji+
7mi6H0FFZ9kxcbiHApxoTd5GUAc5PQtkhsgP+BMofpo7oPWutnHH6GMO4yHTg/BylCL2N4n2nLqA
QbbKn5VtFxQuCOJCXskaCy4GW4t/zGi0nBHVKlVrzto3avHNgMgKNfYDQlJA8opJIs1fCb/irkuK
chPwxwFddloaphi2448DKeLmfM4q9harb2qRrfUehYa98J8acj4ajyMkignqwwkLVCYyuW2U5QfH
aKm5jp68heI9bN+G95/JTZ8w4J1GuCtXVVnGBfcPFNo7BbvbOAZbvkd+Lsj7u7GvZjHG14SmDkem
1aUr7soIMioy7IJocwzklg03sE81UaL3QULRbkVt+vKn2/knACub5lie/x5tclMMuCXzOmIYUQpr
xAgkUwzAcyabBgTySwhQrmapjuJW71+5emjMEEKCCzGF8My2XRETG0kEhOsLCmIhwRMfpz4CW/dF
ALtnKf34Ilrk7xDIWb6tGMTEmNLhVdwTBk3VQ9ogMy/YAufbmhlwcMY1nY2WXELThhR31vqp5C5p
T+kXhkZpxQiRKJfBkaIoxuPrsEt83P8EUBwGLCYJaOgwevCcU4R0Dd4oASE01Cn4eB9hPgginbwL
QbQ/g/R81GcVoQDsjnID4it4FSCMA92e8ZwjUiKC+bqYW2bwktU6fMhi9bNP/A8r25AKZ/GLGSZI
yDciw0m5KembUHOHJ22ozEz0p3CVWl+HOX+GakoWKRyucJzwFYfX1Hk0iD7k1uLlQiS0nxgk0A/e
DXwurQjVGUQ2SZbgQc6OFWuFxyeH+H6bouNrLcD6oGyPhPwO727Z+m7NALOdnudldaRu8SDReTyz
M/l0NkZn65HHGPLsIHm1xsR5RSqZQPlUjwFTrzxst4a6Q5kA1NE6FMv4TVbfJtj5waLP93sHrrhA
fRLDmCcpaDxnT5Es0t7PNUCx5papSloEU1v45fUuUyVpZI02SewhRKpO9VFfZQUauco9lUtcp5uo
OAmyMPV8fC2+EHOF31CwRPJLa+Pcm23L+kJXJ0bEBMU2SO55yFw3AlpPqaXcWIusiH/zcY9TGdtm
kzA1De+C77zU0qxHVS+PisURPyiVBVJrvbofOyjTTPp0NKUseSzxZZfCu44QW4x9I4mATMqtls8q
PW4haIRw1h/T0acyrVVL1XVtHrwgpeiosyfmz3ZLJt0cAZ7Bf16X/C1gjZMy6zzLYO8Cadx4Talt
5zX/JbqNPYjPcvNRDTvzBf9iMa6QEJBgrPjQ7XnuHJghNi8y9Ed1AZVAkpHWt1l9/pj/PBylXHyv
TR1qSpMvo256/IUCwdpwq0zKbyD1z0UIt+g1Dge8E12B4UJMEuDfSbDOOZ56HjOAVFIEiFy1ggmH
17DXJGW10H4mHpgGDOqCJLqP327Pg/cnm8iHCyG+qRMS5V/RLGO0SGpQWyL3N2V77msaYYS/06MQ
djEMRM0p69VQcAKZgdQALzcXukvHj8DKLh74sz3nZae/LUwsFAJnJ2qSp4S6WhwVEbhKNGkP34Lo
vRRuOwPHGHbuK9n9KX3XpKU3OUUX8ewgdPwdEDPhU6mWxFOWesomePGCR6J1+H1J/rgB8LQvFcdB
NbxEPQCCprBooy5Kkd7L1pkugI9m07img9egFhHZytRy1UsZ5bBaiVto103dY8NyyChjGfZ6B3OI
jpSjjoGKx6W2aNGtKb4+hd8QY3BZFC4+IHq9F+bM6QaaVCMtUKRszK1jiOP/4Dedkdc6xYDWUpud
ns7DaybHthFAOnD9dOs8NQK1+/OeTc5rndb8w7PtB9Lkv3hbxnFlFQ1gEvj+xmWgbHTblYtyOBxG
rgSnnyUy0Z0z9jlGhuJukYCqNnl7lBN3UYiBxPYXgA+h3Fy6pdOFTd2ML5vqilNaXxiPp3XqIXgr
guOgovzZbZmT2gGG6n+ADi29DmevNQTqyqRM49s5tZzUMQbXzQC/bB4a5LDd7F0XqDcGhSXBQQvG
v7rj3sL5oePn05ZALFeAKe9Yr+dkHd9uDiK/NECW2PJExso/Zl88BNF5J1lydN7yjnjvGlnb0JIi
fVpGBQUoDePuOOv7EsQJOPxWl/Tr27vPzX2ZdMCVOyu7f6I06cwT9faeOoW1BmHxFi4PGUz1KgVh
hiYt9Ow3yHcbFaOZ8y8YpyB2sTMVP/KtDPWQTR4L+By5Wrg4r0kYjUpVImGfuZdEKb5OpuExOVQ7
snfW5lXH2/76wwijyCMsaIIXL+5qNkrAWppYNIltWwm9ELfzSJ5vr5tfr8FDxtPJ0v/SI74uRq6+
CYTHexESzwqxuppf4OnbHnVD9jtM2LeDU2HEllBYg6Sq+8BrsKQYQQUFo1hIqoUNoD679oYIxCVB
eqDQ0LM7QTdH+vzNUqKuh9RsvnTzUpxi0yhfUXPqzuCxXouPKbH7PyN97MA9Jceq/WcuW1Ps5+cA
xIB2zk8Ewh3lMlppuV0bL1ge6iuOuG/cU8MknVMhW41k650hINh0H0soUQP15NWvkzhmk3vD8Vr1
Ezxr+QNEuMfsNznQOTVKB8Pmc2mTYZrCAjBTN0xzWY4S68/N0EPhL/R8Ddg5xWzHVDMQRbOp0Ych
W1MlsswEHnvIzk0AmvqJXBoVU72seHYWZ7s1MWuqGs7rtK8TED04edHoAYAzt0LYKt2p/DB5Q7x7
kEhJg5TsA7ABsl5xyJmp1o2xdqQx8LB+wTlzojS8v36RM7Bggsyc6ZCkfSW2xrN0DUun8H76ECh4
FCOPohCAXBbw19NmYARKFqqVvCUm0gUTRJg4AQythdkf+D3UnjFsxtQ9uCB86yJCO98A8cP/5STR
vYpdx91MmlZBeXLHoU5qa08ZKqeUPrAfjvoq+gzPpnrUJMb7Wn4UCpyFnbmJznV555aVZ0i97NnA
5OAEyq8oHlZJILrE58WIsMci+3ArZ2UR8+GupBtpY7PZOMdV39+7CJdNj2rrNZo6SXebpTIQeov6
F41cG/bEEF4WFYUTfv1/4eYmHs3tC8WW1KdRhQtXmkC0LPeB/wK2mHv7giwFaPAF9RmpkNDlbhEV
wcgjxw4gs9hGOFdxlBk0OQpHIODiOxHSZlM8g4z67LJ/czbM/PInc3je9xr9uBTcPyowg/FT3bBM
JTRBeyXDBm2FqvCAT7NNBWWw81rhr+5Mkxbk4psiWn5sXpWL5KRPt4bG0mnasXbhBg/wwTSB0dIu
dAjNCVMwFj2yawLRr3OBTO2ZAek2BTvlJA0hL5/4j3fFZ2coze7IR/VokVTLl+22KSs2UP1rhP/D
o8LwFMfX0tfU19kn2B2GaQsgw1oP/ARdg7tb7K43Pz83bldz4/4jX6DpuyyT0xMOHPonDT9Xng7b
++61SBOwIjqzAHsV7t19u8HzIR6XfjeTxHb7h2WVsbvZ4mIEP7NZ5sZiKxBOqRhri+XTsPpSj5qS
4axU8rFe9scbOm/iXIeDlhKPYWGHXni2h9SxWAqrDlWRFpyYXvbP55U3eNvB5Tgk33rX2ZKim2RP
nSZRzC/AaEvhDJbrsMGJE5Fgf/An31GXw9TlhhvHSUVnBRQfEvQcUs9QS9PP3DlPf6eCO2UXcy1w
35xeWLL/HZO3fnqU+yVo1MA52hwmkYyAH2zkk1cslT81aHD6TQp1LExNNIc7/IoYiZqFofy7XFa9
YG5/fIy1FGwPb/Pnn8xjnnp0pSxtVWy2116HaJybBY+TUw7zhAg/3p6Zoxa/hjmrB0EdoJHq/Tyc
4awxRbmx/HqcvoKz09bTxdWDgPHkU5AQzrgVnCMRElfIVEGEpu6BrR25GMNRwedeZIqKADetR13n
NvSn6654GV/zRGEQf3pXiwDXaIOBlFyx4XhTwO5qfuQEwcxo+FRhTy9FoOY47AZnHlZYAfObQTJj
u7cW5ztNwp+nf/xqnylEa+tiUaPZUUpMWQ3Nb5NzUD/Fp/Wewh/a0yTr7Ab4bTvDwJKJlqeH6b1b
xrel9PxyNxY8QPQ0gISDOg77p91QWIekINxuQelbyNQfB4g8cJzcmpAuvAt0RVcEmwnU1hpVeZFV
f142mv0LLyJIl2hHF3j/DwxCAxT02guXigkO8CpQ9QLBRlXuiPuq0moRSdIIM7bEMatfFs+AlsAh
yOkT5P+LvpS9p5px/ul6Pad0/4UbUAOyb+XMEL9HM5VPRPzG2sfhjsdLhIXjvGeucMr3ZCn07bBU
Nf3yHpr1CGOzvCIZv7TW4Wc6+/Hlkrjk8NKZaSytVZCF2GW+TMqFS3tglWi0GzRC+t65G4Co8cES
onGKNxAwdRRjChUmT77ENMB6BeXoRyI7QMT4WQnAiyECmWZNgFtkz0lb3HbhQvnp67xQS6UScSDh
FWlE2IALpPQaINDhAxbC4ubm/gvjAaQpykSGzoje/03PrYBLFwoJSOsHu6H6xxHHMFbxMQ7UwV2q
rZyepi0GrKRG+q9wq3D3oL1sY2ACCmh2qPB/ou6ojnBlS6xFcUqZmYYaPkjb5V4FikKSg+F18gAu
WqvyuwArCrBFRcRI0/+v//8bWVTusZqUyRT86U1o1AozbKxpgLSgmK1+YrKNDKPUUGlYV+0Fq2ao
Q9YrY5kKJO3YIZT+pZPHls2i6WVb4UYwH8BJiwdkiX5CMa3pQRv8SyO/eqE2BEyT/fU1GY2hdCU5
CGjqUCJeJ19DakHYSmsrUuZBcM08LsYfK1pkTh1XiHLa9h+ePtDC4mulek69IklBBxxGLTJLRbgJ
ZhPpfWlKBWhkr5+e7ioPNz8qy7LT+H/803MqezxIgQKxKjhfc7aDIEh4LrqlZuAWg7JK1Be3m1K2
0DVGcNpfickLuRVJv6bhVWbcjgTd5i+A0GdRsfePL2A2Bv0gdV2/x7Ws4oA2Y69vZ+9EEHWB7BKS
5kEFgQ1wI1GsttEO/AYECYmpPVbtwaMZ23HGiLcPqE/c4VZcgEqkiu4R+ZX151FJ6wlv8QBMYenw
eWHn48Qa1Q/wRFeZn8jjeoYnXx709RLgvoXre0ygvIedcjzjoT5NgNZFY6z4Qg7QnsbJ6kRhKOCg
geW9KJrFlGxlmszxw+ciX+hCMCwXWNw5Q8mBNRmEDO58QfHH7VOgSOCmHcbK60NuWIM+IHCK0c6A
RYL31VYcfJBwFEzgbJ4wYi1eePd6AAJ9EhrH+ChEcejYKKLYG0UC9dgvcs4nPENsXNyitLTXvpld
CKIv9LLZa/AvXr63Vim5sgnzuGdoWK41Rd8JF3rmP6KtgnyhOZ7E+NMseHSoI0iArw1hS0p16pyI
T5BaH/ycvqfDDUAgQT2RvWlmPlCiJlMP4ulYPgQ3xscTBzfv4EmW6q3VlfktgDlChBqncp5X5c21
y89ywjOw++JVznk/rKa3Jqei3E3s3ljNyiHql4ltFU1NOJ3qkBpMEPopt+k2CT7b7ecCavJBzj1w
H1d+jusTxBBhjkNY1k4Sor3ZDeTc8/+Uxx7mRYjIfJ07HwRUheIWW2kATssFx0WMfeN876JceQMX
GfHqgDAeDlcseZbdxVekrl60+LiPB/rgsmuAbzrxREPn0A5HQceEV5UHYZCpo+c7GveED2UzdBHp
ZZlAUOgGyiwX+Iv5xIQ4awyEI38kGzjWvhGewVq/pLQTy/H1lDxUp5M24DMceFLTbn0lWxjDG9Jf
O9miabYixGMbmPuSnlkzalrhV1dN880lra1OdLV3C3Vw2LnWDjJ5CkPfn2pYn9K9JbNcp4zlDscl
aUC2eoXZSVa11sQyPWbbTAIRyAcY29C7fc4SILm+TbKruziMMsuEzaw1/rF1pojmGRORqxQvOopP
6nDBa7/1ziZOBY9ODSN5OKpfMNC3+lmANESzQuJ9xvDHcxqWksTJoVG94hAQpObJekbQBX8fzRwz
9OhuLHmCJmomabNh0bNkp8KHhc1HDTYXwAKcTh5e2oBpBXvJAiDWwrVMGZtydHudaqg7gG198zb2
EHcgPhGsX/wpeHkSuNzkVpaqsUZAonybgCIMB3qrI5NbMii/rsWmU5uFHuIaTG/KdoEUdxRYJ4az
MBzZzEyyMY+V3zitdwTqIwFSLp9PADJUOr9PQIweILCsmNWt3Tue5CQ73mlSNz4VJ2wCFSFIspZr
by7UGbqu0ZrFaR+Bw4E0PqwZNt/E172coNN17r8ib3y3x6VhMXHm1RhS3ti0NGQtdEzGlPhxR1bc
OphyGKU3ql7mQXMY9Dx6pWp9wK+m8krDRsJEBR5RcXMhU/Mt6uRgf/eXNvfCoeonJlA3G9go25CX
FnV1okPpuTokIsozD3CRE5V9ALVZvt1fWuOerBh6TNTk9kNE5dLXaffd7YUOmXTypH1LruZr5Vae
rFZllFsXHefH2Ap7nP9N2+/+/Zeln7swSFfwN3eis2cJak/JcIJ5pryAMo7iwzGGmyPmKGiy58Ji
jyrAcXM54jde3GdwcWJnymvm1od9ehXyyyzmiUXfqBpxbjOjwSNv7GkVzIDLxx3DhaIQ/fDqeCwG
skFcvmBqwUdajqM6CNKydvHNdDLD23mcLBsO8o+lUDiSmBG5fJ4lJOOb8G9WV/G3G2N6iU9QH1+t
Vh3kYC6Bud8dHf41Ih4UfpbjmL/9ZMuHzW3hFZvFEtX+vsiWAT/96Fitjn0u8a0sYtqiTDiI/6VK
KqHYWxrY2dk+WJV2vk2wcCL29r6UNI1oXd3qbLz3/97EzWAfGNchqUwljjM25tMuwwQ8AOQonrv1
SZcTqDSvCLlwaXNpJif/wO6vwdFHNGDO93CDA3rj3U4oOwaudoMsgQ+JwaYdmOblS6Qfho4lVC+O
HELeCwlSRCbdoQZGskwoIxfvAwnWFFSv6vhE/WKnxiGwTJYzhBCyyipEWAOgImd9ma8sm9nKDr/b
o2vNid/BkX8WW8vaAFqFucbtkHz6SghjISdSdUgwG+nA3Ov6mlvl5x4TMlxUaMmdnZOE6woYFmce
Fsyuvf+EIQVRXtsRLUOKrpZonCo4hseVayToTj4q+Ik/6zrhiHf5V3SyBH0wDlMxWIBx+R0ZPeAb
DuMuq4EtvLBbGvpR59A5vUkALxpI52If8VPGFwl2bCfl+enpCfKKBaB5YaiLBaLLFYMxBgFvl+Jf
7X1IOqjp7WtMcUWXz7H6rC5o//0Upbxnfa1hjms1q4MXasPbfKZiX4/0PnjRe3eQudwR87h/+c0W
jHuUpGR1Pr54rYfBxy553Rf89+rU16yKYfGMzRphVZ+eHEK6f3FRuFKq1Lb3sYzoPAegy9Unnktl
i8EgK+eLJVDRZm3ZdGynZ/eAkBLxHbxCDDNQhNxZinquYUVX6gB76lqF4cNTZ+kC39SD2L5YYVv4
jmGjmRCTt9xJGGCfSa9nc3QolMNsT7X4XMR/IVZbDtF37d1ehFPGPcR60pa6Rojr5rxC2H1aFOui
fn0TxKhVHPyNb/BO3X5Cc6yylRgmnrLzEgWfZVymJWaAR6K/hUJnFd3CnodlQSEWM8jQQCsvK1JU
WM6Lw6RMO86HFgWWsuzTHxbevKKNGUmP3km08XVSGANwDP5/EYHFmzBNlhSZ8tqFkdhmXRgZOeI5
EUJndBoyxIQbrh0sqGNtLjDnKLdAK/FBEQM+F/h/0bRgOq40vpfG/gFaIC4Mjax85DLvARxCy8Nr
SCugU9yIx+2WV7ed7XsyGrAf1HhH++kIaQLosN7L+NbBerxvFpu07A5u1oEe0uCjwfqcVCmoZxcv
+C8NzkMyPSKhDMRL/xK6B0l4EbywJuHJF2jBXAyqiXRFgCzgOR5523rURTdAvmp8Eo6q3S5zbrgo
lJq4DMXl46Edwd3rDSDwuADB9ptqTvbUeoZBL+29uyD1JXqaY24Uuy2veNbZ6RGSJGPB/DZgO5HA
+7LCTa6xDezmo0LfDqHqR0y0IEQXxhCoozLz6OVKQ0HA+CP/gQFhiooj0m0+wKJRjBdaxGQ3DJDV
48l2d8CW+0Xt6moFsGEbj+qs7q8TOXBy9I1YrlBXRFB/zrfrkwouIwUH/8OvSsm1Lkbpq0aYoLsX
8i1oulliwAiqZv9GA+JutesTLacfjDMQmmVtwqE4Df9KhVSyeOTKOnujSx70ayJDgH4pM1cwNcNj
fW2eN6BO5irDL9n0vWJzlH3mUAIS9VXDqWpOBgUeRHhjxkj8a2G+kwDJxe0OWoDkwCHudEdC/qJI
kuFvmaknfR4rCZW2f2ia5ElMWvqbvGhMxaiDDFw6P5pfgCOxNwkl68mYFycCOZWqHsV2AcXkFpfg
1BAdiXpCjCiOS8aXExdv0CcZL6vKDkUB4dKQ8nTXHqJaAUKqY7lq6h70QNk6u4/cY4Ov+VVvBaiU
a8bnJVFC0vGXVpzVEdIxJKagP38H2uUF6gearO9DtXg5W6KrcuEAp8QXa+EuBrbgnAtgZxnjNbJ3
DAY8Nbz+sLVitZq0eecA1t39oRpU0UM3QU5RoDj+lxF6aMCBJB94kx2WQiczFLfVlAMpgQXJkDkz
NfWxdmYsLT6GR+GZpA60j7kuASz2fGucg9J7+5eh7FLFrD2I1Oy71+CDzyjsdeLTNNkEOh55D0yD
aTmEwbAJocPVAj1k65JBhwbLO/rvM4zMxlTAM7YMU00PhpAKL2AvbKYk6t9tHJdVl6UOoZuavmPf
8WskqczI9QXOFyS9OCOa4d4FLY+NPbIzkO5PRoRideSfJRp6dzt5wfYaST2hraB+AT2Jr4J9MnEH
8ozsliWBwFoZwm0BH7Bxr/xLgL2AjlyXgUFgoLzL0syyUI6EROmBGvLhJxSJLqPhC1hIrZ9+JNhc
XYpiWFbM8vUdBZ8HWxWSlGDzDeK0pre/E47OuU11bmJvwEuR9AtwgEtcEnKrMNRop94inTyTlXQc
tOGhkOO2ilO7v/R7T/cLZ+fQBfIgtXH36qEWXBIHw39+ewR2aE1HKpkeojMpXKO3a11EbON6tsV5
CsVdZmmHB/Vyvu5UYJwWA5qO+8Vcp3vrrPA+b/i2a6XoEjO7hJKLTgbd/t4tuVjs6ftJza9aX6V7
OnQ6fNtBvhYrDJqe5xM70GxCdvJnnwtU5O/iWakuk51nfhEOPYrV9z4uJuQ4BzFCuZvi12pXhXI7
Soskndfo4hmtOcSZgtr74G3aLYYEQifI3zfvaspV7Tqa3GuBIwLHlvaDgx/f8U9JgcKyk7VZy1Z0
UaA6hnF7BfjI7dhYSOboV2Yb8PCFFjQhp0DplOwoD+wV1iuf62Kd74AdUJ38QqOL7IeFNiXaYowo
S6pzBfSk6PS1uSj4Dk5ZUUVcf5afSjXTQZQwWmYveoQJI8GL2hNQ3vBJiKh32EIpw4APRXoXNrKr
kS8kfsFx2kt+CGea9JTlr5ZZPInDIRsmy+Vk+34a/PCmg2ZYNPgs2cKUDOPzkyyWCfTMjBR9H91e
KQnr/DWV2hO9YOYUYdzilfyUhRpXyOMkhsHY6ddGRtMBLFUMc76mIJ44kovGOhIP6cFZU0rGnsbx
Ktz0aO6/opgtMNbgfj8Q4BcvxrwG3alSmV+bhtiTXZ58cnImsjzf1ebNNs58HorhEJ6I8Sv+1HGC
xAAoX1HvavwZUa90uVEYN341aFrwwZRfi8NELLXRio2GheiMjUkRm7j4P8XG3Mbzv91L1UlaYcLj
ztpaX9Uguolm6EyVU3wz5LTlTCWV7/uY+s7MFfJTwm5LYZuaOCbPyPfnla3kRVXYBZxsO25PG3lc
ioureBtHmPUSMunZ0uO7Dm8U6Wqg5Sn0JAs253Zh3HQFgJfYbFgWOXGGrko6hVLZwIViLf6gKwgw
L00AavEUNuReRQH6+OoleJ8nhqMERtwdJBglDvi2D9LZfZm4jU0QfRNnQ4xUJMHNwyKn/Cc5uyIM
qPrXeFGNedb9wBvoL8iYz7VvRShhKTwx2+Ioyfa6pAa2D3vkQ0vZZeW/o3f5YwstISeCL6ZXO1gh
DDzyRDMTOxNFoH2CJHtPivDxHekNgA1cbFpcV7GJuemttR5gpykt8pX39v8sy8GLktjYkWtLlMEI
J/3JTPUmdOzBHUWV9Gw9m6nJPWRM1xrewTiYb0wLG8J9U7y1yVh0mSSFDQI5wriMaHWPpZV17Fbl
cCYsi1KnhfneDwWZpart2kfAPnLnCKaQhfEiYN7ocOZTzitRMzGy7/swazTAc1Z58Gr8RuqJOLee
i4Yfhrt/gKBxE79eH9v7iRMxUtDqAaqbrIMZZStj9eq6CoYtSZhCmCyKwnkNi9Cimrp8NST0ChUB
flG3W19tEplp0EorMEiMEhbNPHmjb28yLKhmHbdF6rsD2M8v3UeeXmDvqlJUe9NQmirBHWbkPN+Q
DwKWtIeLErZhRW+vMwwUUHaXsBIZBlH3p2Nx6nlHGX1Jk7pDb5MpTYCKn2ESCsgApw/vsiBLug2B
lftnxI3C74C5b8hLnIeX5EYR3vArdyi2cVjNdLDEQVMIkrh1RKyDlSgcsk/j2JaRYuCRcJOiZbVE
+FxBewVjpYwP/FW9/xrVUuylt0p0nYfvFdMlfCkFrtSFhoV5EtCsTgFNvtsMDkP3bouEkAFRlifq
g049EFy+vvX0gxPXzNKKsOYD2KOiktcXfQT0hsREV2oR8seRuRC/NlTo42Zq7P5+pBkUZVEb6nWO
VC0X9NS4rMf4pEdyMtChExM3M3NlUSKJoNqYVpZTkdJK68IPc69lgiV3ra9yTLtuQn8FYJytFFvt
5YL8whRZkc+eSBuWkGgBfvq7hSYcVDQp7x8RbziEi649ikdBajXSTRMEg8c/jyDdQXKKIkx8QpnE
lXWNnWxuBsbsRMb6T5c7b72U8qt3kt/6c61WdbHywcx4eeE6sXHv74Qlk2vcUo7bB4JuzFk9jdOz
3azLxOUxVLgWSwwcghFAq0Sy9tiFZwo6zCOF+lKCH5PtjeSuCRHuezkLmWgxIGtO5o3Cj8/c2DZk
cdkDdRgASuPB2ySPtQzd8v7A4XXD9YFzFKheb1WcUgOdtWibyrl73Dm/GJjRqa66md3Li7c4ZR5z
JapX7SATY8eZUgYCnSpJxyfqm0y78GgrOhsepH2M/q/RGzp3BIMmIQ+s9mUUPkWk6QZ16Vgtd4yu
b8qq2U2k3tj4v7hJGvn60zFc8o89nPbVkxbXlNJ2l2NX
`pragma protect end_protected

